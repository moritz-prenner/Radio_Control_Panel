PK
     Y�#\rB�. .    cirkitFile.json{"raven_core_version":15,"hardware_version":0,"pin_to_graph":{"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_0":["pin-type-component_23fc18c5-afdf-44c6-a2e0-9396684812ec_0"],"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_1":["pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_0"],"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_2":["pin-type-component_50742c29-992b-4903-90b0-2b0e050f33c3_0","pin-type-component_f2a462ab-ea50-4a2a-b82c-f46be08c644d_0"],"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_3":[],"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_4":[],"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_5":[],"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_6":[],"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_7":[],"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_8":["pin-type-component_50742c29-992b-4903-90b0-2b0e050f33c3_3"],"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_9":["pin-type-component_50742c29-992b-4903-90b0-2b0e050f33c3_4"],"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_10":["pin-type-component_50742c29-992b-4903-90b0-2b0e050f33c3_1"],"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_11":["pin-type-component_f2a462ab-ea50-4a2a-b82c-f46be08c644d_1"],"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_12":[],"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_13":[],"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_14":[],"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_15":["pin-type-component_f2a462ab-ea50-4a2a-b82c-f46be08c644d_4"],"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_16":["pin-type-component_f2a462ab-ea50-4a2a-b82c-f46be08c644d_3"],"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_17":["pin-type-component_a445ac75-2887-4038-8380-8331f88b6ecf_1","pin-type-component_bcb0cdc5-b2e5-4225-bf8a-97ffe0688c08_1"],"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_18":["pin-type-component_a445ac75-2887-4038-8380-8331f88b6ecf_0"],"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_19":["pin-type-component_bcb0cdc5-b2e5-4225-bf8a-97ffe0688c08_0"],"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_20":["pin-type-component_12231b65-3028-489c-8193-bed54f57003c_0"],"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_21":["pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_0"],"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_22":[],"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_23":["pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_2","pin-type-component_12231b65-3028-489c-8193-bed54f57003c_2","pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_2"],"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_24":["pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_1","pin-type-component_12231b65-3028-489c-8193-bed54f57003c_1","pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_1"],"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_25":[],"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_26":[],"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_27":[],"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_28":[],"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_29":[],"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_30":[],"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_31":[],"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_32":[],"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_33":[],"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_34":[],"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_35":[],"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_36":[],"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_37":["pin-type-component_23fc18c5-afdf-44c6-a2e0-9396684812ec_1","pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_3","pin-type-component_12231b65-3028-489c-8193-bed54f57003c_3","pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_3"],"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_38":[],"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_39":["pin-type-component_99487ac9-98f3-4f19-a8d0-ef91c7362ee4_1","pin-type-component_438418ac-e5ac-420c-b686-a2307c39075f_0","pin-type-component_e45d07ab-a776-4a31-8726-2d647a05518a_0"],"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_40":[],"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_41":[],"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_42":[],"pin-type-component_12231b65-3028-489c-8193-bed54f57003c_0":["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_20"],"pin-type-component_12231b65-3028-489c-8193-bed54f57003c_1":["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_24"],"pin-type-component_12231b65-3028-489c-8193-bed54f57003c_2":["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_23"],"pin-type-component_12231b65-3028-489c-8193-bed54f57003c_3":["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_37"],"pin-type-component_12231b65-3028-489c-8193-bed54f57003c_4":["pin-type-component_438418ac-e5ac-420c-b686-a2307c39075f_1"],"pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_0":["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_21"],"pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_1":["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_24"],"pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_2":["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_23"],"pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_3":["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_37"],"pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_4":["pin-type-component_e45d07ab-a776-4a31-8726-2d647a05518a_1"],"pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_0":["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_1"],"pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_1":["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_24"],"pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_2":["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_23"],"pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_3":["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_37"],"pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_4":["pin-type-component_99487ac9-98f3-4f19-a8d0-ef91c7362ee4_0"],"pin-type-component_a445ac75-2887-4038-8380-8331f88b6ecf_0":["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_18"],"pin-type-component_a445ac75-2887-4038-8380-8331f88b6ecf_1":["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_17"],"pin-type-component_bcb0cdc5-b2e5-4225-bf8a-97ffe0688c08_0":["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_19"],"pin-type-component_bcb0cdc5-b2e5-4225-bf8a-97ffe0688c08_1":["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_17"],"pin-type-component_f2a462ab-ea50-4a2a-b82c-f46be08c644d_0":["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_2"],"pin-type-component_f2a462ab-ea50-4a2a-b82c-f46be08c644d_1":["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_11"],"pin-type-component_f2a462ab-ea50-4a2a-b82c-f46be08c644d_2":[],"pin-type-component_f2a462ab-ea50-4a2a-b82c-f46be08c644d_3":["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_16"],"pin-type-component_f2a462ab-ea50-4a2a-b82c-f46be08c644d_4":["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_15"],"pin-type-component_50742c29-992b-4903-90b0-2b0e050f33c3_0":["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_2"],"pin-type-component_50742c29-992b-4903-90b0-2b0e050f33c3_1":["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_10"],"pin-type-component_50742c29-992b-4903-90b0-2b0e050f33c3_2":[],"pin-type-component_50742c29-992b-4903-90b0-2b0e050f33c3_3":["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_8"],"pin-type-component_50742c29-992b-4903-90b0-2b0e050f33c3_4":["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_9"],"pin-type-component_23fc18c5-afdf-44c6-a2e0-9396684812ec_0":["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_0"],"pin-type-component_23fc18c5-afdf-44c6-a2e0-9396684812ec_1":["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_37"],"pin-type-component_99487ac9-98f3-4f19-a8d0-ef91c7362ee4_0":["pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_4"],"pin-type-component_99487ac9-98f3-4f19-a8d0-ef91c7362ee4_1":["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_39"],"pin-type-component_438418ac-e5ac-420c-b686-a2307c39075f_0":["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_39"],"pin-type-component_438418ac-e5ac-420c-b686-a2307c39075f_1":["pin-type-component_12231b65-3028-489c-8193-bed54f57003c_4"],"pin-type-component_e45d07ab-a776-4a31-8726-2d647a05518a_0":["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_39"],"pin-type-component_e45d07ab-a776-4a31-8726-2d647a05518a_1":["pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_4"]},"pin_to_color":{"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_0":"#010067","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_1":"#95003A","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_2":"#007DB5","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_3":"#000000","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_4":"#000000","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_5":"#000000","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_6":"#000000","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_7":"#000000","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_8":"#683D3B","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_9":"#FF029D","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_10":"#5FAD4E","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_11":"#008F9C","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_12":"#000000","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_13":"#000000","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_14":"#000000","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_15":"#968AE8","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_16":"#FF74A3","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_17":"#6A826C","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_18":"#00AE7E","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_19":"#C28C9F","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_20":"#FF937E","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_21":"#001544","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_22":"#000000","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_23":"#FFE502","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_24":"#91D0CB","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_25":"#000000","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_26":"#000000","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_27":"#000000","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_28":"#000000","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_29":"#000000","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_30":"#000000","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_31":"#000000","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_32":"#000000","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_33":"#000000","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_34":"#000000","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_35":"#000000","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_36":"#000000","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_37":"#9E008E","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_38":"#000000","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_39":"#A75740","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_40":"#000000","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_41":"#000000","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_42":"#000000","pin-type-component_12231b65-3028-489c-8193-bed54f57003c_0":"#FF937E","pin-type-component_12231b65-3028-489c-8193-bed54f57003c_1":"#91D0CB","pin-type-component_12231b65-3028-489c-8193-bed54f57003c_2":"#FFE502","pin-type-component_12231b65-3028-489c-8193-bed54f57003c_3":"#9E008E","pin-type-component_12231b65-3028-489c-8193-bed54f57003c_4":"#01FFFE","pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_0":"#001544","pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_1":"#91D0CB","pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_2":"#FFE502","pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_3":"#9E008E","pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_4":"#FE8900","pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_0":"#95003A","pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_1":"#91D0CB","pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_2":"#FFE502","pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_3":"#9E008E","pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_4":"#98FF52","pin-type-component_a445ac75-2887-4038-8380-8331f88b6ecf_0":"#00AE7E","pin-type-component_a445ac75-2887-4038-8380-8331f88b6ecf_1":"#6A826C","pin-type-component_bcb0cdc5-b2e5-4225-bf8a-97ffe0688c08_0":"#C28C9F","pin-type-component_bcb0cdc5-b2e5-4225-bf8a-97ffe0688c08_1":"#6A826C","pin-type-component_f2a462ab-ea50-4a2a-b82c-f46be08c644d_0":"#007DB5","pin-type-component_f2a462ab-ea50-4a2a-b82c-f46be08c644d_1":"#008F9C","pin-type-component_f2a462ab-ea50-4a2a-b82c-f46be08c644d_2":"#000000","pin-type-component_f2a462ab-ea50-4a2a-b82c-f46be08c644d_3":"#FF74A3","pin-type-component_f2a462ab-ea50-4a2a-b82c-f46be08c644d_4":"#968AE8","pin-type-component_50742c29-992b-4903-90b0-2b0e050f33c3_0":"#007DB5","pin-type-component_50742c29-992b-4903-90b0-2b0e050f33c3_1":"#5FAD4E","pin-type-component_50742c29-992b-4903-90b0-2b0e050f33c3_2":"#000000","pin-type-component_50742c29-992b-4903-90b0-2b0e050f33c3_3":"#683D3B","pin-type-component_50742c29-992b-4903-90b0-2b0e050f33c3_4":"#FF029D","pin-type-component_23fc18c5-afdf-44c6-a2e0-9396684812ec_0":"#010067","pin-type-component_23fc18c5-afdf-44c6-a2e0-9396684812ec_1":"#9E008E","pin-type-component_99487ac9-98f3-4f19-a8d0-ef91c7362ee4_0":"#98FF52","pin-type-component_99487ac9-98f3-4f19-a8d0-ef91c7362ee4_1":"#A75740","pin-type-component_438418ac-e5ac-420c-b686-a2307c39075f_0":"#A75740","pin-type-component_438418ac-e5ac-420c-b686-a2307c39075f_1":"#01FFFE","pin-type-component_e45d07ab-a776-4a31-8726-2d647a05518a_0":"#A75740","pin-type-component_e45d07ab-a776-4a31-8726-2d647a05518a_1":"#FE8900"},"pin_to_state":{"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_0":"neutral","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_1":"neutral","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_2":"neutral","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_3":"neutral","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_4":"neutral","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_5":"neutral","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_6":"neutral","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_7":"neutral","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_8":"neutral","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_9":"neutral","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_10":"neutral","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_11":"neutral","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_12":"neutral","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_13":"neutral","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_14":"neutral","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_15":"neutral","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_16":"neutral","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_17":"neutral","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_18":"neutral","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_19":"neutral","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_20":"neutral","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_21":"neutral","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_22":"neutral","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_23":"neutral","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_24":"neutral","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_25":"neutral","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_26":"neutral","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_27":"neutral","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_28":"neutral","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_29":"neutral","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_30":"neutral","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_31":"neutral","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_32":"neutral","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_33":"neutral","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_34":"neutral","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_35":"neutral","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_36":"neutral","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_37":"neutral","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_38":"neutral","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_39":"neutral","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_40":"neutral","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_41":"neutral","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_42":"neutral","pin-type-component_12231b65-3028-489c-8193-bed54f57003c_0":"neutral","pin-type-component_12231b65-3028-489c-8193-bed54f57003c_1":"neutral","pin-type-component_12231b65-3028-489c-8193-bed54f57003c_2":"neutral","pin-type-component_12231b65-3028-489c-8193-bed54f57003c_3":"neutral","pin-type-component_12231b65-3028-489c-8193-bed54f57003c_4":"neutral","pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_0":"neutral","pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_1":"neutral","pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_2":"neutral","pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_3":"neutral","pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_4":"neutral","pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_0":"neutral","pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_1":"neutral","pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_2":"neutral","pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_3":"neutral","pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_4":"neutral","pin-type-component_a445ac75-2887-4038-8380-8331f88b6ecf_0":"neutral","pin-type-component_a445ac75-2887-4038-8380-8331f88b6ecf_1":"neutral","pin-type-component_bcb0cdc5-b2e5-4225-bf8a-97ffe0688c08_0":"neutral","pin-type-component_bcb0cdc5-b2e5-4225-bf8a-97ffe0688c08_1":"neutral","pin-type-component_f2a462ab-ea50-4a2a-b82c-f46be08c644d_0":"neutral","pin-type-component_f2a462ab-ea50-4a2a-b82c-f46be08c644d_1":"neutral","pin-type-component_f2a462ab-ea50-4a2a-b82c-f46be08c644d_2":"neutral","pin-type-component_f2a462ab-ea50-4a2a-b82c-f46be08c644d_3":"neutral","pin-type-component_f2a462ab-ea50-4a2a-b82c-f46be08c644d_4":"neutral","pin-type-component_50742c29-992b-4903-90b0-2b0e050f33c3_0":"neutral","pin-type-component_50742c29-992b-4903-90b0-2b0e050f33c3_1":"neutral","pin-type-component_50742c29-992b-4903-90b0-2b0e050f33c3_2":"neutral","pin-type-component_50742c29-992b-4903-90b0-2b0e050f33c3_3":"neutral","pin-type-component_50742c29-992b-4903-90b0-2b0e050f33c3_4":"neutral","pin-type-component_23fc18c5-afdf-44c6-a2e0-9396684812ec_0":"neutral","pin-type-component_23fc18c5-afdf-44c6-a2e0-9396684812ec_1":"neutral","pin-type-component_99487ac9-98f3-4f19-a8d0-ef91c7362ee4_0":"neutral","pin-type-component_99487ac9-98f3-4f19-a8d0-ef91c7362ee4_1":"neutral","pin-type-component_438418ac-e5ac-420c-b686-a2307c39075f_0":"neutral","pin-type-component_438418ac-e5ac-420c-b686-a2307c39075f_1":"neutral","pin-type-component_e45d07ab-a776-4a31-8726-2d647a05518a_0":"neutral","pin-type-component_e45d07ab-a776-4a31-8726-2d647a05518a_1":"neutral"},"next_color_idx":23,"wires_placed_in_order":[["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_0","pin-type-component_23fc18c5-afdf-44c6-a2e0-9396684812ec_0"],["pin-type-component_23fc18c5-afdf-44c6-a2e0-9396684812ec_1","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_37"],["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_37","pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_3"],["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_37","pin-type-component_12231b65-3028-489c-8193-bed54f57003c_3"],["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_37","pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_3"],["pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_1","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_33"],["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_33","pin-type-component_12231b65-3028-489c-8193-bed54f57003c_1"],["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_33","pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_1"],["pin-type-component_12231b65-3028-489c-8193-bed54f57003c_2","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_31"],["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_31","pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_2"],["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_31","pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_2"],["pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_4","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_39"],["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_39","pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_4"],["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_39","pin-type-component_12231b65-3028-489c-8193-bed54f57003c_4"],["pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_0","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_1"],["pin-type-component_12231b65-3028-489c-8193-bed54f57003c_0","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_20"],["pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_0","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_21"],["pin-type-component_12231b65-3028-489c-8193-bed54f57003c_2","pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_2"],["pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_2","pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_2"],["pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_2","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_23"],["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_23","pin-type-component_12231b65-3028-489c-8193-bed54f57003c_2"],["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_23","pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_2"],["pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_1","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_24"],["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_24","pin-type-component_12231b65-3028-489c-8193-bed54f57003c_1"],["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_24","pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_1"],["pin-type-component_50742c29-992b-4903-90b0-2b0e050f33c3_0","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_2"],["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_2","pin-type-component_f2a462ab-ea50-4a2a-b82c-f46be08c644d_0"],["pin-type-component_a445ac75-2887-4038-8380-8331f88b6ecf_1","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_17"],["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_17","pin-type-component_bcb0cdc5-b2e5-4225-bf8a-97ffe0688c08_1"],["pin-type-component_a445ac75-2887-4038-8380-8331f88b6ecf_0","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_18"],["pin-type-component_bcb0cdc5-b2e5-4225-bf8a-97ffe0688c08_0","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_19"],["pin-type-component_f2a462ab-ea50-4a2a-b82c-f46be08c644d_1","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_11"],["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_10","pin-type-component_50742c29-992b-4903-90b0-2b0e050f33c3_1"],["pin-type-component_50742c29-992b-4903-90b0-2b0e050f33c3_4","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_9"],["pin-type-component_50742c29-992b-4903-90b0-2b0e050f33c3_3","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_8"],["pin-type-component_f2a462ab-ea50-4a2a-b82c-f46be08c644d_3","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_16"],["pin-type-component_f2a462ab-ea50-4a2a-b82c-f46be08c644d_4","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_15"],["pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_4","pin-type-component_99487ac9-98f3-4f19-a8d0-ef91c7362ee4_0"],["pin-type-component_99487ac9-98f3-4f19-a8d0-ef91c7362ee4_1","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_39"],["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_39","pin-type-component_438418ac-e5ac-420c-b686-a2307c39075f_0"],["pin-type-component_438418ac-e5ac-420c-b686-a2307c39075f_1","pin-type-component_12231b65-3028-489c-8193-bed54f57003c_4"],["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_39","pin-type-component_e45d07ab-a776-4a31-8726-2d647a05518a_0"],["pin-type-component_e45d07ab-a776-4a31-8726-2d647a05518a_1","pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_4"]],"wires_removed_and_placed_in_order":[[[],[["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_0","pin-type-component_23fc18c5-afdf-44c6-a2e0-9396684812ec_0"]]],[[],[["pin-type-component_23fc18c5-afdf-44c6-a2e0-9396684812ec_1","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_37"]]],[[],[["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_37","pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_3"]]],[[],[["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_37","pin-type-component_12231b65-3028-489c-8193-bed54f57003c_3"]]],[[],[["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_37","pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_3"]]],[[],[["pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_1","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_33"]]],[[],[["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_33","pin-type-component_12231b65-3028-489c-8193-bed54f57003c_1"]]],[[],[["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_33","pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_1"]]],[[],[["pin-type-component_12231b65-3028-489c-8193-bed54f57003c_2","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_31"]]],[[],[["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_31","pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_2"]]],[[],[["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_31","pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_2"]]],[[],[["pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_4","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_39"]]],[[],[["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_39","pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_4"]]],[[],[["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_39","pin-type-component_12231b65-3028-489c-8193-bed54f57003c_4"]]],[[],[["pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_0","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_1"]]],[[],[["pin-type-component_12231b65-3028-489c-8193-bed54f57003c_0","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_20"]]],[[],[["pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_0","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_21"]]],[[["pin-type-component_12231b65-3028-489c-8193-bed54f57003c_2","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_31"],["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_31","pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_2"],["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_31","pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_2"]],[["pin-type-component_12231b65-3028-489c-8193-bed54f57003c_2","pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_2"],["pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_2","pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_2"]]],[[],[["pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_2","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_23"]]],[[["pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_2","pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_2"]],[]],[[["pin-type-component_12231b65-3028-489c-8193-bed54f57003c_2","pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_2"]],[]],[[],[["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_23","pin-type-component_12231b65-3028-489c-8193-bed54f57003c_2"]]],[[],[["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_23","pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_2"]]],[[["pin-type-component_12231b65-3028-489c-8193-bed54f57003c_1","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_33"]],[]],[[["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_33","pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_1"]],[]],[[["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_33","pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_1"]],[]],[[],[["pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_1","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_24"]]],[[],[["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_24","pin-type-component_12231b65-3028-489c-8193-bed54f57003c_1"]]],[[],[["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_24","pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_1"]]],[[],[["pin-type-component_50742c29-992b-4903-90b0-2b0e050f33c3_0","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_2"]]],[[],[["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_2","pin-type-component_f2a462ab-ea50-4a2a-b82c-f46be08c644d_0"]]],[[],[["pin-type-component_a445ac75-2887-4038-8380-8331f88b6ecf_1","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_17"]]],[[],[["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_17","pin-type-component_bcb0cdc5-b2e5-4225-bf8a-97ffe0688c08_1"]]],[[],[["pin-type-component_a445ac75-2887-4038-8380-8331f88b6ecf_0","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_18"]]],[[],[["pin-type-component_bcb0cdc5-b2e5-4225-bf8a-97ffe0688c08_0","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_19"]]],[[],[["pin-type-component_f2a462ab-ea50-4a2a-b82c-f46be08c644d_1","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_11"]]],[[],[["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_10","pin-type-component_50742c29-992b-4903-90b0-2b0e050f33c3_1"]]],[[],[["pin-type-component_50742c29-992b-4903-90b0-2b0e050f33c3_4","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_9"]]],[[],[["pin-type-component_50742c29-992b-4903-90b0-2b0e050f33c3_3","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_8"]]],[[],[["pin-type-component_f2a462ab-ea50-4a2a-b82c-f46be08c644d_3","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_16"]]],[[],[["pin-type-component_f2a462ab-ea50-4a2a-b82c-f46be08c644d_4","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_15"]]],[[["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_39","pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_4"]],[]],[[["pin-type-component_12231b65-3028-489c-8193-bed54f57003c_4","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_39"]],[]],[[["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_39","pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_4"]],[]],[[],[["pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_4","pin-type-component_99487ac9-98f3-4f19-a8d0-ef91c7362ee4_0"]]],[[],[["pin-type-component_99487ac9-98f3-4f19-a8d0-ef91c7362ee4_1","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_39"]]],[[],[["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_39","pin-type-component_438418ac-e5ac-420c-b686-a2307c39075f_0"]]],[[],[["pin-type-component_438418ac-e5ac-420c-b686-a2307c39075f_1","pin-type-component_12231b65-3028-489c-8193-bed54f57003c_4"]]],[[],[["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_39","pin-type-component_e45d07ab-a776-4a31-8726-2d647a05518a_0"]]],[[],[["pin-type-component_e45d07ab-a776-4a31-8726-2d647a05518a_1","pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_4"]]]],"arduino_state":"arduino_off","pin_to_uid":{"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_0":"0000000000000000","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_1":"0000000000000005","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_2":"0000000000000008","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_3":"_","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_4":"_","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_5":"_","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_6":"_","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_7":"_","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_8":"0000000000000015","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_9":"0000000000000014","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_10":"0000000000000013","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_11":"0000000000000012","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_12":"_","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_13":"_","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_14":"_","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_15":"0000000000000017","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_16":"0000000000000016","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_17":"0000000000000009","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_18":"0000000000000010","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_19":"0000000000000011","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_20":"0000000000000006","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_21":"0000000000000007","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_22":"_","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_23":"0000000000000003","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_24":"0000000000000002","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_25":"_","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_26":"_","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_27":"_","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_28":"_","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_29":"_","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_30":"_","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_31":"_","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_32":"_","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_33":"_","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_34":"_","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_35":"_","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_36":"_","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_37":"0000000000000001","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_38":"_","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_39":"0000000000000018","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_40":"_","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_41":"_","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_42":"_","pin-type-component_12231b65-3028-489c-8193-bed54f57003c_0":"0000000000000006","pin-type-component_12231b65-3028-489c-8193-bed54f57003c_1":"0000000000000002","pin-type-component_12231b65-3028-489c-8193-bed54f57003c_2":"0000000000000003","pin-type-component_12231b65-3028-489c-8193-bed54f57003c_3":"0000000000000001","pin-type-component_12231b65-3028-489c-8193-bed54f57003c_4":"0000000000000019","pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_0":"0000000000000007","pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_1":"0000000000000002","pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_2":"0000000000000003","pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_3":"0000000000000001","pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_4":"0000000000000020","pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_0":"0000000000000005","pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_1":"0000000000000002","pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_2":"0000000000000003","pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_3":"0000000000000001","pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_4":"0000000000000004","pin-type-component_a445ac75-2887-4038-8380-8331f88b6ecf_0":"0000000000000010","pin-type-component_a445ac75-2887-4038-8380-8331f88b6ecf_1":"0000000000000009","pin-type-component_bcb0cdc5-b2e5-4225-bf8a-97ffe0688c08_0":"0000000000000011","pin-type-component_bcb0cdc5-b2e5-4225-bf8a-97ffe0688c08_1":"0000000000000009","pin-type-component_f2a462ab-ea50-4a2a-b82c-f46be08c644d_0":"0000000000000008","pin-type-component_f2a462ab-ea50-4a2a-b82c-f46be08c644d_1":"0000000000000012","pin-type-component_f2a462ab-ea50-4a2a-b82c-f46be08c644d_2":"_","pin-type-component_f2a462ab-ea50-4a2a-b82c-f46be08c644d_3":"0000000000000016","pin-type-component_f2a462ab-ea50-4a2a-b82c-f46be08c644d_4":"0000000000000017","pin-type-component_50742c29-992b-4903-90b0-2b0e050f33c3_0":"0000000000000008","pin-type-component_50742c29-992b-4903-90b0-2b0e050f33c3_1":"0000000000000013","pin-type-component_50742c29-992b-4903-90b0-2b0e050f33c3_2":"_","pin-type-component_50742c29-992b-4903-90b0-2b0e050f33c3_3":"0000000000000015","pin-type-component_50742c29-992b-4903-90b0-2b0e050f33c3_4":"0000000000000014","pin-type-component_23fc18c5-afdf-44c6-a2e0-9396684812ec_0":"0000000000000000","pin-type-component_23fc18c5-afdf-44c6-a2e0-9396684812ec_1":"0000000000000001","pin-type-component_99487ac9-98f3-4f19-a8d0-ef91c7362ee4_0":"0000000000000004","pin-type-component_99487ac9-98f3-4f19-a8d0-ef91c7362ee4_1":"0000000000000018","pin-type-component_438418ac-e5ac-420c-b686-a2307c39075f_0":"0000000000000018","pin-type-component_438418ac-e5ac-420c-b686-a2307c39075f_1":"0000000000000019","pin-type-component_e45d07ab-a776-4a31-8726-2d647a05518a_0":"0000000000000018","pin-type-component_e45d07ab-a776-4a31-8726-2d647a05518a_1":"0000000000000020"},"component_id_to_pins":{"91d5d40b-a663-4f86-bb6a-531c98c6974e":["0","1","2","3","4","5","6","7","8","9","10","11","12","13","14","15","16","17","18","19","20","21","22","23","24","25","26","27","28","29","30","31","32","33","34","35","36","37","38","39","40","41","42"],"12231b65-3028-489c-8193-bed54f57003c":["0","1","2","3","4"],"ec8d45f2-93af-4156-af57-a8dad25ff981":["0","1","2","3","4"],"e82ce461-d5a2-4a54-b071-a766699ccc57":["0","1","2","3","4"],"a445ac75-2887-4038-8380-8331f88b6ecf":["0","1"],"bcb0cdc5-b2e5-4225-bf8a-97ffe0688c08":["0","1"],"f2a462ab-ea50-4a2a-b82c-f46be08c644d":["0","1","2","3","4"],"50742c29-992b-4903-90b0-2b0e050f33c3":["0","1","2","3","4"],"23fc18c5-afdf-44c6-a2e0-9396684812ec":["0","1"],"99487ac9-98f3-4f19-a8d0-ef91c7362ee4":["0","1"],"438418ac-e5ac-420c-b686-a2307c39075f":["0","1"],"e45d07ab-a776-4a31-8726-2d647a05518a":["0","1"]},"uid_to_net":{"_":[],"0000000000000000":["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_0","pin-type-component_23fc18c5-afdf-44c6-a2e0-9396684812ec_0"],"0000000000000001":["pin-type-component_12231b65-3028-489c-8193-bed54f57003c_3","pin-type-component_23fc18c5-afdf-44c6-a2e0-9396684812ec_1","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_37","pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_3","pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_3"],"0000000000000003":["pin-type-component_12231b65-3028-489c-8193-bed54f57003c_2","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_23","pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_2","pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_2"],"0000000000000005":["pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_0","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_1"],"0000000000000006":["pin-type-component_12231b65-3028-489c-8193-bed54f57003c_0","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_20"],"0000000000000007":["pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_0","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_21"],"0000000000000002":["pin-type-component_12231b65-3028-489c-8193-bed54f57003c_1","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_24","pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_1","pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_1"],"0000000000000008":["pin-type-component_50742c29-992b-4903-90b0-2b0e050f33c3_0","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_2","pin-type-component_f2a462ab-ea50-4a2a-b82c-f46be08c644d_0"],"0000000000000009":["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_17","pin-type-component_a445ac75-2887-4038-8380-8331f88b6ecf_1","pin-type-component_bcb0cdc5-b2e5-4225-bf8a-97ffe0688c08_1"],"0000000000000010":["pin-type-component_a445ac75-2887-4038-8380-8331f88b6ecf_0","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_18"],"0000000000000011":["pin-type-component_bcb0cdc5-b2e5-4225-bf8a-97ffe0688c08_0","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_19"],"0000000000000012":["pin-type-component_f2a462ab-ea50-4a2a-b82c-f46be08c644d_1","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_11"],"0000000000000013":["pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_10","pin-type-component_50742c29-992b-4903-90b0-2b0e050f33c3_1"],"0000000000000014":["pin-type-component_50742c29-992b-4903-90b0-2b0e050f33c3_4","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_9"],"0000000000000015":["pin-type-component_50742c29-992b-4903-90b0-2b0e050f33c3_3","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_8"],"0000000000000016":["pin-type-component_f2a462ab-ea50-4a2a-b82c-f46be08c644d_3","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_16"],"0000000000000017":["pin-type-component_f2a462ab-ea50-4a2a-b82c-f46be08c644d_4","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_15"],"0000000000000004":["pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_4","pin-type-component_99487ac9-98f3-4f19-a8d0-ef91c7362ee4_0"],"0000000000000018":["pin-type-component_438418ac-e5ac-420c-b686-a2307c39075f_0","pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_39","pin-type-component_99487ac9-98f3-4f19-a8d0-ef91c7362ee4_1","pin-type-component_e45d07ab-a776-4a31-8726-2d647a05518a_0"],"0000000000000019":["pin-type-component_438418ac-e5ac-420c-b686-a2307c39075f_1","pin-type-component_12231b65-3028-489c-8193-bed54f57003c_4"],"0000000000000020":["pin-type-component_e45d07ab-a776-4a31-8726-2d647a05518a_1","pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_4"]},"uid_to_text_label":{"0000000000000000":"Net 0","0000000000000001":"Net 1","0000000000000003":"Net 3","0000000000000005":"Net 5","0000000000000006":"Net 6","0000000000000007":"Net 7","0000000000000002":"Net 2","0000000000000008":"Net 8","0000000000000009":"Net 9","0000000000000010":"Net 10","0000000000000011":"Net 11","0000000000000012":"Net 12","0000000000000013":"Net 13","0000000000000014":"Net 14","0000000000000015":"Net 15","0000000000000016":"Net 16","0000000000000017":"Net 17","0000000000000004":"Net 4","0000000000000018":"Net 18","0000000000000019":"Net 19","0000000000000020":"Net 20"},"all_breadboard_info_list":[],"breadboard_info_list":[],"componentsData":[{"compProperties":{},"position":[610.89295,276.61258999999995],"typeId":"a075aea4-de2b-28dc-4d34-388439862a7a","componentVersion":34,"instanceId":"91d5d40b-a663-4f86-bb6a-531c98c6974e","orientation":"up","circleData":[[557.5,139.99999999999997],[557.5,155.00899999999993],[557.5,170.00899999999993],[557.5,185.00899999999993],[557.5,200.00899999999993],[557.5,215.00899999999993],[557.5,230.00899999999993],[557.5,245.00899999999993],[557.4340000000001,260.0089999999999],[557.4340000000001,275.00899999999996],[557.4340000000001,290.00899999999996],[557.4340000000001,305.00899999999996],[557.4340000000001,320.00899999999996],[557.4340000000001,335.00899999999996],[557.4340000000001,350.00899999999996],[557.4340000000001,365.00899999999996],[557.4340000000001,380.00899999999996],[557.4340000000001,395.00899999999996],[557.4340000000001,410.00899999999996],[557.4340000000001,425.00899999999996],[662.4340000000001,425.00899999999996],[662.4340000000001,410.00899999999996],[662.4340000000001,395.00899999999996],[662.4340000000001,380.00899999999996],[662.4340000000001,365.00899999999996],[662.4340000000001,350.00899999999996],[662.4340000000001,335.00899999999996],[662.4340000000001,320.00899999999996],[662.4340000000001,305.00899999999996],[662.4340000000001,290.00899999999996],[662.4340000000001,275.00899999999996],[662.4340000000001,260.0089999999999],[662.4340000000001,245.00899999999993],[662.4340000000001,230.00899999999993],[662.4340000000001,215.00899999999993],[662.4340000000001,200.00899999999993],[662.4340000000001,185.00899999999993],[662.4340000000001,170.00899999999993],[662.4340000000001,155.00899999999993],[662.4340000000001,140.00899999999993],[594.9343735,425.00938849999994],[609.9343735,425.00938849999994],[624.9343765,425.00938849999994]],"code":"517,folder,{\"name\":\"sketch\",\"id\":\"5b18efba-42ce-4848-9377-7bdd2f9df882\",\"explorerHtmlId\":\"0d0caf7f-5415-4d96-8243-7e74e5947103\",\"nameHtmlId\":\"8444dbbb-5acf-4eca-bb90-e77a8dad3e2e\",\"nameInputHtmlId\":\"9d4dac52-f16f-4cf2-bf64-4d5b3ce8a2ca\",\"explorerChildHtmlId\":\"f4190374-3896-4583-8b43-0a34def375b8\",\"explorerCarrotOpenHtmlId\":\"88c79196-7bec-49a4-8244-8b8c6de3fa14\",\"explorerCarrotClosedHtmlId\":\"82947504-d2fb-41db-ab81-e048d3188ba7\",\"arduinoBoardFqbn\":\"rp2040:rp2040:rpipico\",\"arduinoBoardName\":\"\",\"arduinoPortAddress\":\"\"},2,381,file,{\"name\":\"sketch.ino\",\"id\":\"fbaa1c04-3c15-4868-a2ad-3ec59fc635e8\",\"explorerHtmlId\":\"7d3ae622-88a8-4c9c-b7c2-899ddacd0ad3\",\"nameHtmlId\":\"c32e0592-57cd-4616-8afd-8358eda40155\",\"nameInputHtmlId\":\"72ccdc5a-34c8-4a7d-af25-c27b2583daae\",\"code\":\"void setup() {\\n  // put your setup code here, to run once:\\n\\n}\\n\\nvoid loop() {\\n  // put your main code here, to run repeatedly:\\n\\n}\"},0,252,file,{\"name\":\"documentation.txt\",\"id\":\"172df276-dc73-4104-9d11-c4f86ef778c4\",\"explorerHtmlId\":\"3b6e0319-c245-4e32-9767-cb62cc889ea9\",\"nameHtmlId\":\"1bfb1553-d1eb-4538-9d07-19e16d918f6c\",\"nameInputHtmlId\":\"7ededbe1-781d-450f-81a0-62660725fc6d\",\"code\":\"\"},0,","codeLabelPosition":[610.89295,120.09096499999998],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[915.1004005,185.526839],"typeId":"aae483c6-3d50-4df0-8aab-097e662db2ce","componentVersion":1,"instanceId":"12231b65-3028-489c-8193-bed54f57003c","orientation":"up","circleData":[[872.5,155],[873.649,170.79650000000004],[871.255,189.464],[873.169,207.17449999999997],[872.6904999999999,223.928]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[915.1004005,335.526839],"typeId":"aae483c6-3d50-4df0-8aab-097e662db2ce","componentVersion":1,"instanceId":"ec8d45f2-93af-4156-af57-a8dad25ff981","orientation":"up","circleData":[[872.5,305],[873.649,320.79650000000004],[871.255,339.464],[873.169,357.17449999999997],[872.6904999999999,373.928]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[915.1004005,20.526838999999974],"typeId":"aae483c6-3d50-4df0-8aab-097e662db2ce","componentVersion":1,"instanceId":"e82ce461-d5a2-4a54-b071-a766699ccc57","orientation":"up","circleData":[[872.5,-10.000000000000007],[873.6489999999999,5.79650000000003],[871.2550000000001,24.463999999999988],[873.1689999999999,42.17449999999996],[872.6904999999999,58.92799999999992]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[403.8845244999999,538.012523],"typeId":"481439cd-69fa-4157-bae3-cbd35387bdef","componentVersion":1,"instanceId":"a445ac75-2887-4038-8380-8331f88b6ecf","orientation":"up","circleData":[[377.5,545],[420.27549999999985,545.9105000000001]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[403.8845245000001,628.012523],"typeId":"481439cd-69fa-4157-bae3-cbd35387bdef","componentVersion":1,"instanceId":"bcb0cdc5-b2e5-4225-bf8a-97ffe0688c08","orientation":"up","circleData":[[377.5,635],[420.2755,635.9105000000001]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[378.1786809999999,353.8697840000001],"typeId":"73eff55f-a5c6-450f-b7e9-078fea8511d1","componentVersion":1,"instanceId":"f2a462ab-ea50-4a2a-b82c-f46be08c644d","orientation":"up","circleData":[[407.5,365],[407.5,341.8722439999999],[349.68061,353.43612199999995],[349.68061,330.308366],[351.9933849999999,376.56387800000005]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[378.17868100000004,218.86978399999998],"typeId":"73eff55f-a5c6-450f-b7e9-078fea8511d1","componentVersion":1,"instanceId":"50742c29-992b-4903-90b0-2b0e050f33c3","orientation":"up","circleData":[[407.5,230.00000000000003],[407.5,206.8722439999999],[349.68060999999994,218.43612199999995],[349.68060999999994,195.30836599999998],[351.9933849999998,241.56387800000007]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[422.6067475,-17.174718999999982],"typeId":"115f87dd-3a9c-47f0-b7ba-2c17fa02ee85","componentVersion":1,"instanceId":"23fc18c5-afdf-44c6-a2e0-9396684812ec","orientation":"up","circleData":[[347.5,-9.999999999999993],[497.50000000000017,-9.999999999999993]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Capacitance":{"version":2,"id":"Capacitance","label":"Capacitance","description":"","units":"F","type":"decimal","value":"0.0000001","displayFormat":"input","showOnComp":true,"isVisibleToUser":true}},"position":[1030.012,16.379750000000026],"typeId":"2c229afa-5375-44c6-9069-3781267c16db","componentVersion":1,"instanceId":"99487ac9-98f3-4f19-a8d0-ef91c7362ee4","orientation":"up","circleData":[[1022.5,65],[1037.5345,65]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Capacitance":{"version":2,"id":"Capacitance","label":"Capacitance","description":"","units":"F","type":"decimal","value":"0.0000001","displayFormat":"input","showOnComp":true,"isVisibleToUser":true,"name":"Capacitance","unit":"F","required":true}},"position":[1075.012,46.37974999999996],"typeId":"2c229afa-5375-44c6-9069-3781267c16db","componentVersion":1,"instanceId":"438418ac-e5ac-420c-b686-a2307c39075f","orientation":"up","circleData":[[1067.5,94.99999999999997],[1082.5345,94.99999999999997]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Capacitance":{"version":2,"id":"Capacitance","label":"Capacitance","description":"","units":"F","type":"decimal","value":"0.0000001","displayFormat":"input","showOnComp":true,"isVisibleToUser":true,"name":"Capacitance","unit":"F","required":true}},"position":[1135.012,31.37975000000023],"typeId":"2c229afa-5375-44c6-9069-3781267c16db","componentVersion":1,"instanceId":"e45d07ab-a776-4a31-8726-2d647a05518a","orientation":"up","circleData":[[1127.5,80.00000000000003],[1142.5345,80.00000000000003]],"cirkitStudioVersion":"1.3.3"}],"bounds":{"top":"-51.07444","left":"333.50000","width":"825.63900","height":"723.64577","x":"333.50000","y":"-51.07444"},"cachedBreadboardPrettyViewWires":["{\"color\":\"#010067\",\"startPinId\":\"pin-type-component_23fc18c5-afdf-44c6-a2e0-9396684812ec_0\",\"endPinId\":\"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_0\",\"rawStartPinId\":\"pin-type-component_23fc18c5-afdf-44c6-a2e0-9396684812ec_0\",\"rawEndPinId\":\"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"347.5000000000_-10.0000000000\\\",\\\"332.5000000000_-10.0000000000\\\",\\\"332.5000000000_140.0000000000\\\",\\\"557.5000000000_140.0000000000\\\"]}\"}","{\"color\":\"#9E008E\",\"startPinId\":\"pin-type-component_23fc18c5-afdf-44c6-a2e0-9396684812ec_1\",\"endPinId\":\"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_37\",\"rawStartPinId\":\"pin-type-component_23fc18c5-afdf-44c6-a2e0-9396684812ec_1\",\"rawEndPinId\":\"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_37\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"497.5000000000_-10.0000000000\\\",\\\"707.5000000000_-10.0000000000\\\",\\\"707.5000000000_170.0090000000\\\",\\\"662.4340000000_170.0090000000\\\"]}\"}","{\"color\":\"#9E008E\",\"startPinId\":\"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_37\",\"endPinId\":\"pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_3\",\"rawStartPinId\":\"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_37\",\"rawEndPinId\":\"pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"662.4340000000_170.0090000000\\\",\\\"782.5000000000_170.0090000000\\\",\\\"782.5000000000_42.1745000000\\\",\\\"873.1690000000_42.1745000000\\\"]}\"}","{\"color\":\"#9E008E\",\"startPinId\":\"pin-type-component_12231b65-3028-489c-8193-bed54f57003c_3\",\"endPinId\":\"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_37\",\"rawStartPinId\":\"pin-type-component_12231b65-3028-489c-8193-bed54f57003c_3\",\"rawEndPinId\":\"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_37\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"873.1690000000_207.1745000000\\\",\\\"782.5000000000_207.1745000000\\\",\\\"782.5000000000_170.0090000000\\\",\\\"662.4340000000_170.0090000000\\\"]}\"}","{\"color\":\"#9E008E\",\"startPinId\":\"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_37\",\"endPinId\":\"pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_3\",\"rawStartPinId\":\"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_37\",\"rawEndPinId\":\"pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"662.4340000000_170.0090000000\\\",\\\"782.5000000000_170.0090000000\\\",\\\"782.5000000000_357.1745000000\\\",\\\"873.1690000000_357.1745000000\\\"]}\"}","{\"color\":\"#95003A\",\"startPinId\":\"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_1\",\"endPinId\":\"pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_0\",\"rawStartPinId\":\"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_1\",\"rawEndPinId\":\"pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"557.5000000000_155.0090000000\\\",\\\"527.5000000000_155.0090000000\\\",\\\"527.5000000000_-55.0000000000\\\",\\\"872.5000000000_-55.0000000000\\\",\\\"872.5000000000_-10.0000000000\\\"]}\"}","{\"color\":\"#FF937E\",\"startPinId\":\"pin-type-component_12231b65-3028-489c-8193-bed54f57003c_0\",\"endPinId\":\"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_20\",\"rawStartPinId\":\"pin-type-component_12231b65-3028-489c-8193-bed54f57003c_0\",\"rawEndPinId\":\"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_20\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"872.5000000000_155.0000000000\\\",\\\"1052.5000000000_155.0000000000\\\",\\\"1052.5000000000_455.0000000000\\\",\\\"662.4340000000_455.0000000000\\\",\\\"662.4340000000_425.0090000000\\\"]}\"}","{\"color\":\"#001544\",\"startPinId\":\"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_21\",\"endPinId\":\"pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_0\",\"rawStartPinId\":\"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_21\",\"rawEndPinId\":\"pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"662.4340000000_410.0090000000\\\",\\\"835.0000000000_410.0090000000\\\",\\\"835.0000000000_305.0000000000\\\",\\\"872.5000000000_305.0000000000\\\"]}\"}","{\"color\":\"#FFE502\",\"startPinId\":\"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_23\",\"endPinId\":\"pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_2\",\"rawStartPinId\":\"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_23\",\"rawEndPinId\":\"pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"662.4340000000_380.0090000000\\\",\\\"730.0000000000_380.0090000000\\\",\\\"730.0000000000_24.4640000000\\\",\\\"871.2550000000_24.4640000000\\\"]}\"}","{\"color\":\"#FFE502\",\"startPinId\":\"pin-type-component_12231b65-3028-489c-8193-bed54f57003c_2\",\"endPinId\":\"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_23\",\"rawStartPinId\":\"pin-type-component_12231b65-3028-489c-8193-bed54f57003c_2\",\"rawEndPinId\":\"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_23\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"871.2550000000_189.4640000000\\\",\\\"730.0000000000_189.4640000000\\\",\\\"730.0000000000_380.0090000000\\\",\\\"662.4340000000_380.0090000000\\\"]}\"}","{\"color\":\"#FFE502\",\"startPinId\":\"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_23\",\"endPinId\":\"pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_2\",\"rawStartPinId\":\"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_23\",\"rawEndPinId\":\"pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"662.4340000000_380.0090000000\\\",\\\"730.0000000000_380.0090000000\\\",\\\"730.0000000000_339.4640000000\\\",\\\"871.2550000000_339.4640000000\\\"]}\"}","{\"color\":\"#91D0CB\",\"startPinId\":\"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_24\",\"endPinId\":\"pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_1\",\"rawStartPinId\":\"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_24\",\"rawEndPinId\":\"pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"662.4340000000_365.0090000000\\\",\\\"752.5000000000_365.0090000000\\\",\\\"752.5000000000_5.7965000000\\\",\\\"873.6490000000_5.7965000000\\\"]}\"}","{\"color\":\"#91D0CB\",\"startPinId\":\"pin-type-component_12231b65-3028-489c-8193-bed54f57003c_1\",\"endPinId\":\"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_24\",\"rawStartPinId\":\"pin-type-component_12231b65-3028-489c-8193-bed54f57003c_1\",\"rawEndPinId\":\"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_24\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"873.6490000000_170.7965000000\\\",\\\"827.5000000000_170.7965000000\\\",\\\"827.5000000000_245.0000000000\\\",\\\"752.5000000000_245.0000000000\\\",\\\"752.5000000000_365.0090000000\\\",\\\"662.4340000000_365.0090000000\\\"]}\"}","{\"color\":\"#91D0CB\",\"startPinId\":\"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_24\",\"endPinId\":\"pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_1\",\"rawStartPinId\":\"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_24\",\"rawEndPinId\":\"pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"662.4340000000_365.0090000000\\\",\\\"752.5000000000_365.0090000000\\\",\\\"752.5000000000_320.7965000000\\\",\\\"873.6490000000_320.7965000000\\\"]}\"}","{\"color\":\"#007DB5\",\"startPinId\":\"pin-type-component_50742c29-992b-4903-90b0-2b0e050f33c3_0\",\"endPinId\":\"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_2\",\"rawStartPinId\":\"pin-type-component_50742c29-992b-4903-90b0-2b0e050f33c3_0\",\"rawEndPinId\":\"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"407.5000000000_230.0000000000\\\",\\\"482.5000000000_230.0000000000\\\",\\\"482.5000000000_170.0090000000\\\",\\\"557.5000000000_170.0090000000\\\"]}\"}","{\"color\":\"#007DB5\",\"startPinId\":\"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_2\",\"endPinId\":\"pin-type-component_f2a462ab-ea50-4a2a-b82c-f46be08c644d_0\",\"rawStartPinId\":\"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_2\",\"rawEndPinId\":\"pin-type-component_f2a462ab-ea50-4a2a-b82c-f46be08c644d_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"557.5000000000_170.0090000000\\\",\\\"482.5000000000_170.0090000000\\\",\\\"482.5000000000_365.0000000000\\\",\\\"407.5000000000_365.0000000000\\\"]}\"}","{\"color\":\"#6A826C\",\"startPinId\":\"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_17\",\"endPinId\":\"pin-type-component_a445ac75-2887-4038-8380-8331f88b6ecf_1\",\"rawStartPinId\":\"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_17\",\"rawEndPinId\":\"pin-type-component_a445ac75-2887-4038-8380-8331f88b6ecf_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"557.4340000000_395.0090000000\\\",\\\"482.5000000000_395.0090000000\\\",\\\"482.5000000000_545.0000000000\\\",\\\"420.2755000000_545.0000000000\\\",\\\"420.2755000000_545.9105000000\\\"]}\"}","{\"color\":\"#6A826C\",\"startPinId\":\"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_17\",\"endPinId\":\"pin-type-component_bcb0cdc5-b2e5-4225-bf8a-97ffe0688c08_1\",\"rawStartPinId\":\"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_17\",\"rawEndPinId\":\"pin-type-component_bcb0cdc5-b2e5-4225-bf8a-97ffe0688c08_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"557.4340000000_395.0090000000\\\",\\\"482.5000000000_395.0090000000\\\",\\\"482.5000000000_635.0000000000\\\",\\\"420.2755000000_635.0000000000\\\",\\\"420.2755000000_635.9105000000\\\"]}\"}","{\"color\":\"#00AE7E\",\"startPinId\":\"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_18\",\"endPinId\":\"pin-type-component_a445ac75-2887-4038-8380-8331f88b6ecf_0\",\"rawStartPinId\":\"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_18\",\"rawEndPinId\":\"pin-type-component_a445ac75-2887-4038-8380-8331f88b6ecf_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"557.4340000000_410.0090000000\\\",\\\"332.5000000000_410.0090000000\\\",\\\"332.5000000000_545.0000000000\\\",\\\"377.5000000000_545.0000000000\\\"]}\"}","{\"color\":\"#C28C9F\",\"startPinId\":\"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_19\",\"endPinId\":\"pin-type-component_bcb0cdc5-b2e5-4225-bf8a-97ffe0688c08_0\",\"rawStartPinId\":\"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_19\",\"rawEndPinId\":\"pin-type-component_bcb0cdc5-b2e5-4225-bf8a-97ffe0688c08_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"557.4340000000_425.0090000000\\\",\\\"557.4340000000_680.0000000000\\\",\\\"332.5000000000_680.0000000000\\\",\\\"332.5000000000_635.0000000000\\\",\\\"377.5000000000_635.0000000000\\\"]}\"}","{\"color\":\"#008F9C\",\"startPinId\":\"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_11\",\"endPinId\":\"pin-type-component_f2a462ab-ea50-4a2a-b82c-f46be08c644d_1\",\"rawStartPinId\":\"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_11\",\"rawEndPinId\":\"pin-type-component_f2a462ab-ea50-4a2a-b82c-f46be08c644d_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"557.4340000000_305.0090000000\\\",\\\"520.0000000000_305.0090000000\\\",\\\"520.0000000000_341.8722440000\\\",\\\"407.5000000000_341.8722440000\\\"]}\"}","{\"color\":\"#5FAD4E\",\"startPinId\":\"pin-type-component_50742c29-992b-4903-90b0-2b0e050f33c3_1\",\"endPinId\":\"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_10\",\"rawStartPinId\":\"pin-type-component_50742c29-992b-4903-90b0-2b0e050f33c3_1\",\"rawEndPinId\":\"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_10\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"407.5000000000_206.8722440000\\\",\\\"460.0000000000_206.8722440000\\\",\\\"460.0000000000_290.0090000000\\\",\\\"557.4340000000_290.0090000000\\\"]}\"}","{\"color\":\"#FF029D\",\"startPinId\":\"pin-type-component_50742c29-992b-4903-90b0-2b0e050f33c3_4\",\"endPinId\":\"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_9\",\"rawStartPinId\":\"pin-type-component_50742c29-992b-4903-90b0-2b0e050f33c3_4\",\"rawEndPinId\":\"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_9\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"351.9933850000_241.5638780000\\\",\\\"332.5000000000_241.5638780000\\\",\\\"332.5000000000_275.0090000000\\\",\\\"557.4340000000_275.0090000000\\\"]}\"}","{\"color\":\"#683D3B\",\"startPinId\":\"pin-type-component_50742c29-992b-4903-90b0-2b0e050f33c3_3\",\"endPinId\":\"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_8\",\"rawStartPinId\":\"pin-type-component_50742c29-992b-4903-90b0-2b0e050f33c3_3\",\"rawEndPinId\":\"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_8\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"349.6806100000_195.3083660000\\\",\\\"349.6806100000_155.0000000000\\\",\\\"512.5000000000_155.0000000000\\\",\\\"512.5000000000_260.0090000000\\\",\\\"557.4340000000_260.0090000000\\\"]}\"}","{\"color\":\"#FF74A3\",\"startPinId\":\"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_16\",\"endPinId\":\"pin-type-component_f2a462ab-ea50-4a2a-b82c-f46be08c644d_3\",\"rawStartPinId\":\"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_16\",\"rawEndPinId\":\"pin-type-component_f2a462ab-ea50-4a2a-b82c-f46be08c644d_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"557.4340000000_380.0090000000\\\",\\\"452.5000000000_380.0090000000\\\",\\\"452.5000000000_305.0000000000\\\",\\\"332.5000000000_305.0000000000\\\",\\\"332.5000000000_330.3083660000\\\",\\\"349.6806100000_330.3083660000\\\"]}\"}","{\"color\":\"#968AE8\",\"startPinId\":\"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_15\",\"endPinId\":\"pin-type-component_f2a462ab-ea50-4a2a-b82c-f46be08c644d_4\",\"rawStartPinId\":\"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_15\",\"rawEndPinId\":\"pin-type-component_f2a462ab-ea50-4a2a-b82c-f46be08c644d_4\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"557.4340000000_365.0090000000\\\",\\\"512.5000000000_365.0090000000\\\",\\\"512.5000000000_440.0000000000\\\",\\\"302.5000000000_440.0000000000\\\",\\\"302.5000000000_376.5638780000\\\",\\\"351.9933850000_376.5638780000\\\"]}\"}","{\"color\":\"#98FF52\",\"startPinId\":\"pin-type-component_99487ac9-98f3-4f19-a8d0-ef91c7362ee4_0\",\"endPinId\":\"pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_4\",\"rawStartPinId\":\"pin-type-component_99487ac9-98f3-4f19-a8d0-ef91c7362ee4_0\",\"rawEndPinId\":\"pin-type-component_e82ce461-d5a2-4a54-b071-a766699ccc57_4\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1022.5000000000_65.0000000000\\\",\\\"1022.5000000000_72.5000000000\\\",\\\"872.5000000000_72.5000000000\\\",\\\"872.5000000000_65.0000000000\\\",\\\"872.6905000000_65.0000000000\\\",\\\"872.6905000000_58.9280000000\\\"]}\"}","{\"color\":\"#A75740\",\"startPinId\":\"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_39\",\"endPinId\":\"pin-type-component_99487ac9-98f3-4f19-a8d0-ef91c7362ee4_1\",\"rawStartPinId\":\"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_39\",\"rawEndPinId\":\"pin-type-component_99487ac9-98f3-4f19-a8d0-ef91c7362ee4_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"662.4340000000_140.0090000000\\\",\\\"662.4340000000_95.0000000000\\\",\\\"1037.5345000000_95.0000000000\\\",\\\"1037.5345000000_65.0000000000\\\"]}\"}","{\"color\":\"#A75740\",\"startPinId\":\"pin-type-component_438418ac-e5ac-420c-b686-a2307c39075f_0\",\"endPinId\":\"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_39\",\"rawStartPinId\":\"pin-type-component_438418ac-e5ac-420c-b686-a2307c39075f_0\",\"rawEndPinId\":\"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_39\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1067.5000000000_95.0000000000\\\",\\\"662.4340000000_95.0000000000\\\",\\\"662.4340000000_140.0090000000\\\"]}\"}","{\"color\":\"#A75740\",\"startPinId\":\"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_39\",\"endPinId\":\"pin-type-component_e45d07ab-a776-4a31-8726-2d647a05518a_0\",\"rawStartPinId\":\"pin-type-component_91d5d40b-a663-4f86-bb6a-531c98c6974e_39\",\"rawEndPinId\":\"pin-type-component_e45d07ab-a776-4a31-8726-2d647a05518a_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"662.4340000000_140.0090000000\\\",\\\"662.4340000000_95.0000000000\\\",\\\"1037.5000000000_95.0000000000\\\",\\\"1037.5000000000_125.0000000000\\\",\\\"1127.5000000000_125.0000000000\\\",\\\"1127.5000000000_80.0000000000\\\"]}\"}","{\"color\":\"#01FFFE\",\"startPinId\":\"pin-type-component_12231b65-3028-489c-8193-bed54f57003c_4\",\"endPinId\":\"pin-type-component_438418ac-e5ac-420c-b686-a2307c39075f_1\",\"rawStartPinId\":\"pin-type-component_12231b65-3028-489c-8193-bed54f57003c_4\",\"rawEndPinId\":\"pin-type-component_438418ac-e5ac-420c-b686-a2307c39075f_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"872.6905000000_223.9280000000\\\",\\\"842.5000000000_223.9280000000\\\",\\\"842.5000000000_260.0000000000\\\",\\\"1082.5345000000_260.0000000000\\\",\\\"1082.5345000000_95.0000000000\\\"]}\"}","{\"color\":\"#FE8900\",\"startPinId\":\"pin-type-component_e45d07ab-a776-4a31-8726-2d647a05518a_1\",\"endPinId\":\"pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_4\",\"rawStartPinId\":\"pin-type-component_e45d07ab-a776-4a31-8726-2d647a05518a_1\",\"rawEndPinId\":\"pin-type-component_ec8d45f2-93af-4156-af57-a8dad25ff981_4\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1142.5345000000_80.0000000000\\\",\\\"1142.5345000000_477.5000000000\\\",\\\"902.5000000000_477.5000000000\\\",\\\"902.5000000000_373.9280000000\\\",\\\"872.6905000000_373.9280000000\\\"]}\"}"],"projectDescription":""}PK
     Y�#\               jsons/PK
     Y�#\Y��c|7  |7     jsons/user_defined.json{"type":"user_defined","version":"0.0.1","subtypes":[{"subtypeName":"Raspberry Pi Pico","category":["User Defined"],"userDefined":true,"id":"a075aea4-de2b-28dc-4d34-388439862a7a","fqbn":"rp2040:rp2040:rpipico","subtypeDescription":"","subtypePic":"04079d65-5a5d-4b08-9f2d-4934008ae210.png","iconPic":"c73ef27d-6394-4828-a75f-205a980bbd83.png","imageLocation":"local_cache","componentVersion":34,"pinInfo":{"numDisplayCols":"8.26781","numDisplayRows":"20.86955","pins":[{"uniquePinIdString":"0","positionMil":"57.43750,1954.22810","isAnchorPin":true,"label":"GP0"},{"uniquePinIdString":"1","positionMil":"57.43750,1854.16810","isAnchorPin":false,"label":"GP1"},{"uniquePinIdString":"2","positionMil":"57.43750,1754.16810","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"3","positionMil":"57.43750,1654.16810","isAnchorPin":false,"label":"GP2"},{"uniquePinIdString":"4","positionMil":"57.43750,1554.16810","isAnchorPin":false,"label":"GP3"},{"uniquePinIdString":"5","positionMil":"57.43750,1454.16810","isAnchorPin":false,"label":"GP4"},{"uniquePinIdString":"6","positionMil":"57.43750,1354.16810","isAnchorPin":false,"label":"GP5"},{"uniquePinIdString":"7","positionMil":"57.43750,1254.16810","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"8","positionMil":"56.99750,1154.16810","isAnchorPin":false,"label":"GP6"},{"uniquePinIdString":"9","positionMil":"56.99750,1054.16810","isAnchorPin":false,"label":"GP7"},{"uniquePinIdString":"10","positionMil":"56.99750,954.16810","isAnchorPin":false,"label":"GP8"},{"uniquePinIdString":"11","positionMil":"56.99750,854.16810","isAnchorPin":false,"label":"GP9"},{"uniquePinIdString":"12","positionMil":"56.99750,754.16810","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"13","positionMil":"56.99750,654.16810","isAnchorPin":false,"label":"GP10"},{"uniquePinIdString":"14","positionMil":"56.99750,554.16810","isAnchorPin":false,"label":"GP11"},{"uniquePinIdString":"15","positionMil":"56.99750,454.16810","isAnchorPin":false,"label":"GP12"},{"uniquePinIdString":"16","positionMil":"56.99750,354.16810","isAnchorPin":false,"label":"GP13"},{"uniquePinIdString":"17","positionMil":"56.99750,254.16810","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"18","positionMil":"56.99750,154.16810","isAnchorPin":false,"label":"GP14"},{"uniquePinIdString":"19","positionMil":"56.99750,54.16810","isAnchorPin":false,"label":"GP15"},{"uniquePinIdString":"20","positionMil":"756.99750,54.16810","isAnchorPin":false,"label":"GP16"},{"uniquePinIdString":"21","positionMil":"756.99750,154.16810","isAnchorPin":false,"label":"GP17"},{"uniquePinIdString":"22","positionMil":"756.99750,254.16810","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"23","positionMil":"756.99750,354.16810","isAnchorPin":false,"label":"GP18"},{"uniquePinIdString":"24","positionMil":"756.99750,454.16810","isAnchorPin":false,"label":"GP19"},{"uniquePinIdString":"25","positionMil":"756.99750,554.16810","isAnchorPin":false,"label":"GP20"},{"uniquePinIdString":"26","positionMil":"756.99750,654.16810","isAnchorPin":false,"label":"GP21"},{"uniquePinIdString":"27","positionMil":"756.99750,754.16810","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"28","positionMil":"756.99750,854.16810","isAnchorPin":false,"label":"GP22"},{"uniquePinIdString":"29","positionMil":"756.99750,954.16810","isAnchorPin":false,"label":"RUN"},{"uniquePinIdString":"30","positionMil":"756.99750,1054.16810","isAnchorPin":false,"label":"GP26"},{"uniquePinIdString":"31","positionMil":"756.99750,1154.16810","isAnchorPin":false,"label":"GP27"},{"uniquePinIdString":"32","positionMil":"756.99750,1254.16810","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"33","positionMil":"756.99750,1354.16810","isAnchorPin":false,"label":"GP28"},{"uniquePinIdString":"34","positionMil":"756.99750,1454.16810","isAnchorPin":false,"label":"ADC_VREF"},{"uniquePinIdString":"35","positionMil":"756.99750,1554.16810","isAnchorPin":false,"label":"3V3"},{"uniquePinIdString":"36","positionMil":"756.99750,1654.16810","isAnchorPin":false,"label":"3V3_EN"},{"uniquePinIdString":"37","positionMil":"756.99750,1754.16810","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"38","positionMil":"756.99750,1854.16810","isAnchorPin":false,"label":"VSYS"},{"uniquePinIdString":"39","positionMil":"756.99750,1954.16810","isAnchorPin":false,"label":"VBUS"},{"uniquePinIdString":"40","positionMil":"306.99999,54.16551","isAnchorPin":false,"label":"pin 41"},{"uniquePinIdString":"41","positionMil":"406.99999,54.16551","isAnchorPin":false,"label":"pin 42"},{"uniquePinIdString":"42","positionMil":"507.00001,54.16551","isAnchorPin":false,"label":"pin 43"}],"pinType":"wired"},"properties":[],"hasComponentImageSvg":true,"componentImageSvgUrl":"https://abacasstorageaccnt.blob.core.windows.net/cirkit/9eb97c9b-93be-48e5-ab72-785b9faebafd.svg","propertiesV2":[]},{"subtypeName":"seven segment display","category":["User Defined"],"id":"aae483c6-3d50-4df0-8aab-097e662db2ce","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"c3d75dd9-81e0-4ecb-9109-310dbcf70c9d.png","iconPic":"c7f8a6b2-5f4f-47a7-84b3-7bbc451b7ab1.png","hasComponentImageSvg":false,"componentImageSvgUrl":"","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.85172","numDisplayRows":"6.85172","pins":[{"uniquePinIdString":"0","positionMil":"58.58333,546.09826","isAnchorPin":true,"label":"CS"},{"uniquePinIdString":"1","positionMil":"66.24333,440.78826","isAnchorPin":false,"label":"CLK"},{"uniquePinIdString":"2","positionMil":"50.28333,316.33826","isAnchorPin":false,"label":"DIN"},{"uniquePinIdString":"3","positionMil":"63.04333,198.26826","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"4","positionMil":"59.85333,86.57826","isAnchorPin":false,"label":"VCC"}],"pinType":"wired"},"properties":[],"propertiesV2":[]},{"subtypeName":"seven segment display","category":["User Defined"],"id":"aae483c6-3d50-4df0-8aab-097e662db2ce","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"c3d75dd9-81e0-4ecb-9109-310dbcf70c9d.png","iconPic":"c7f8a6b2-5f4f-47a7-84b3-7bbc451b7ab1.png","hasComponentImageSvg":false,"componentImageSvgUrl":"","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.85172","numDisplayRows":"6.85172","pins":[{"uniquePinIdString":"0","positionMil":"58.58333,546.09826","isAnchorPin":true,"label":"CS"},{"uniquePinIdString":"1","positionMil":"66.24333,440.78826","isAnchorPin":false,"label":"CLK"},{"uniquePinIdString":"2","positionMil":"50.28333,316.33826","isAnchorPin":false,"label":"DIN"},{"uniquePinIdString":"3","positionMil":"63.04333,198.26826","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"4","positionMil":"59.85333,86.57826","isAnchorPin":false,"label":"VCC"}],"pinType":"wired"},"properties":[],"propertiesV2":[]},{"subtypeName":"seven segment display","category":["User Defined"],"id":"aae483c6-3d50-4df0-8aab-097e662db2ce","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"c3d75dd9-81e0-4ecb-9109-310dbcf70c9d.png","iconPic":"c7f8a6b2-5f4f-47a7-84b3-7bbc451b7ab1.png","hasComponentImageSvg":false,"componentImageSvgUrl":"","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.85172","numDisplayRows":"6.85172","pins":[{"uniquePinIdString":"0","positionMil":"58.58333,546.09826","isAnchorPin":true,"label":"CS"},{"uniquePinIdString":"1","positionMil":"66.24333,440.78826","isAnchorPin":false,"label":"CLK"},{"uniquePinIdString":"2","positionMil":"50.28333,316.33826","isAnchorPin":false,"label":"DIN"},{"uniquePinIdString":"3","positionMil":"63.04333,198.26826","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"4","positionMil":"59.85333,86.57826","isAnchorPin":false,"label":"VCC"}],"pinType":"wired"},"properties":[],"propertiesV2":[]},{"subtypeName":"push button","category":["User Defined"],"id":"481439cd-69fa-4157-bae3-cbd35387bdef","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"be1ff175-690b-4799-aad0-0ab57f9a01ac.png","iconPic":"a7a20d0b-f771-49dd-a52a-92c84cdc73c6.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.66667","numDisplayRows":"4.60784","pins":[{"uniquePinIdString":"0","positionMil":"157.43667,183.80882","isAnchorPin":true,"label":"pin1"},{"uniquePinIdString":"1","positionMil":"442.60667,177.73882","isAnchorPin":false,"label":"pin2"}],"pinType":"wired"},"properties":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"push button","category":["User Defined"],"id":"481439cd-69fa-4157-bae3-cbd35387bdef","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"be1ff175-690b-4799-aad0-0ab57f9a01ac.png","iconPic":"a7a20d0b-f771-49dd-a52a-92c84cdc73c6.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.66667","numDisplayRows":"4.60784","pins":[{"uniquePinIdString":"0","positionMil":"157.43667,183.80882","isAnchorPin":true,"label":"pin1"},{"uniquePinIdString":"1","positionMil":"442.60667,177.73882","isAnchorPin":false,"label":"pin2"}],"pinType":"wired"},"properties":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"EC11 Rotary Encoder","category":["User Defined"],"id":"73eff55f-a5c6-450f-b7e9-078fea8511d1","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"e7e47810-abf9-4bb0-84d9-bf12c3babd78.png","iconPic":"9eaf56c3-a2ed-4703-8e91-9b98c221ec28.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"4.58627","numDisplayRows":"4.95813","pins":[{"uniquePinIdString":"0","positionMil":"424.78896,173.70506","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"424.78896,327.89010","isAnchorPin":false,"label":"SW"},{"uniquePinIdString":"2","positionMil":"39.32636,250.79758","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"3","positionMil":"39.32636,404.98262","isAnchorPin":false,"label":"DT"},{"uniquePinIdString":"4","positionMil":"54.74486,96.61254","isAnchorPin":false,"label":"CLK"}],"pinType":"wired"},"properties":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"EC11 Rotary Encoder","category":["User Defined"],"id":"73eff55f-a5c6-450f-b7e9-078fea8511d1","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"e7e47810-abf9-4bb0-84d9-bf12c3babd78.png","iconPic":"9eaf56c3-a2ed-4703-8e91-9b98c221ec28.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"4.58627","numDisplayRows":"4.95813","pins":[{"uniquePinIdString":"0","positionMil":"424.78896,173.70506","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"424.78896,327.89010","isAnchorPin":false,"label":"SW"},{"uniquePinIdString":"2","positionMil":"39.32636,250.79758","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"3","positionMil":"39.32636,404.98262","isAnchorPin":false,"label":"DT"},{"uniquePinIdString":"4","positionMil":"54.74486,96.61254","isAnchorPin":false,"label":"CLK"}],"pinType":"wired"},"properties":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"switch_off","category":["User Defined"],"id":"115f87dd-3a9c-47f0-b7ba-2c17fa02ee85","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"5ccbe72c-6fd5-45d2-8118-bee80363f106.png","iconPic":"e4bf1f14-66df-463a-8792-8567b691137d.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"10.06303","numDisplayRows":"3.18663","pins":[{"uniquePinIdString":"0","positionMil":"2.43985,111.50004","isAnchorPin":true,"label":"1"},{"uniquePinIdString":"1","positionMil":"1002.43985,111.50004","isAnchorPin":false,"label":"2"}],"pinType":"wired"},"properties":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Ceramic Capacitor","subtypeDescription":"","id":"2c229afa-5375-44c6-9069-3781267c16db","subtypePic":"7c9bed20-c7d7-43dc-b689-820375f46db8.png","category":["Basic"],"userDefined":false,"pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"44.10000,0.00000","endPositionMil":"44.10000,-200.00000","isAnchorPin":true,"label":"pin0"},{"uniquePinIdString":"1","startPositionMil":"144.33000,0.00000","endPositionMil":"144.33000,-200.00000","isAnchorPin":false,"label":"pin1"}],"numDisplayCols":"1.88360","numDisplayRows":"2.48270","pinType":"movable"},"properties":[{"type":"double","name":"Capacitance","value":"0.0000001","unit":"F","showOnComp":true,"required":true}],"iconPic":"7ade412b-fa94-47ea-987a-d6c9baa14438.png","componentVersion":1,"imageLocation":"local_cache","hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Ceramic Capacitor","subtypeDescription":"","id":"2c229afa-5375-44c6-9069-3781267c16db","subtypePic":"7c9bed20-c7d7-43dc-b689-820375f46db8.png","category":["Basic"],"userDefined":false,"pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"44.10000,0.00000","endPositionMil":"44.10000,-200.00000","isAnchorPin":true,"label":"pin0"},{"uniquePinIdString":"1","startPositionMil":"144.33000,0.00000","endPositionMil":"144.33000,-200.00000","isAnchorPin":false,"label":"pin1"}],"numDisplayCols":"1.88360","numDisplayRows":"2.48270","pinType":"movable"},"properties":[{"type":"double","name":"Capacitance","value":"0.0000001","unit":"F","showOnComp":true,"required":true}],"iconPic":"7ade412b-fa94-47ea-987a-d6c9baa14438.png","componentVersion":1,"imageLocation":"local_cache","hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Ceramic Capacitor","subtypeDescription":"","id":"2c229afa-5375-44c6-9069-3781267c16db","subtypePic":"7c9bed20-c7d7-43dc-b689-820375f46db8.png","category":["Basic"],"userDefined":false,"pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"44.10000,0.00000","endPositionMil":"44.10000,-200.00000","isAnchorPin":true,"label":"pin0"},{"uniquePinIdString":"1","startPositionMil":"144.33000,0.00000","endPositionMil":"144.33000,-200.00000","isAnchorPin":false,"label":"pin1"}],"numDisplayCols":"1.88360","numDisplayRows":"2.48270","pinType":"movable"},"properties":[{"type":"double","name":"Capacitance","value":"0.0000001","unit":"F","showOnComp":true,"required":true}],"iconPic":"7ade412b-fa94-47ea-987a-d6c9baa14438.png","componentVersion":1,"imageLocation":"local_cache","hasComponentImageSvg":false,"componentImageSvgUrl":""}]}PK
     Y�#\               images/PK
     Y�#\��9�� �� /   images/04079d65-5a5d-4b08-9f2d-4934008ae210.png�PNG

   IHDR  �  �   ��R�   	pHYs  \F  \F�CA  ��IDATx���|e� ��%��4�-��.�ʞ2DF�TP�u�D_Sо�
*��nQ�R�,Y*���Y(�h�J���=�x$m�\���~b���i.��=�=����ӧ���D���R Y��Bn�(����I)�����ˀP�����K����!����u��M��j�㧎���&.
�Qן�2 T����-������q⎵��㻦M� !?���*'''��XwpA1A��̀t�ɓ�NHh��l�ݻw�$���0@H��,۲eKӞ={ڝ�p����Z�w2�3-��~�ر�M�4)��8�+J�>��?��S2��X�]I�9o�_���F���(����3�{���m��̉ܜ����J�����Y��t@�O0�#�b�.������'O���=\��\-} �,E'	��ɓ}(	���Kb!?����*���k���8ܖ�srr\v�yEA�C�ɛ5kf��<K1OPp�Qʰp�#L�ȯ(����ߝXvDn��䜛��T�y �T�L%��=���3'N�H��ϡNw��6@ȏ0�#�JHH8p�TN)W��W~��(�����x�e�A��y��AP)�s�ﷸc��8�BQR\R����6L�ȯHG����W�ݱ�eGs5�Ow�� ���e�t��e��x���\�~�Ş˹c���8�?�Z����;��$\���СC�ejYS.�6���;��<y���l��j���(�o��~ ?B~�	��6��-��b��(H�+�Ӂ�2��s�,�H�92IPs��Y���l��3L���,9'sp�����`_g)8IaG>��0���8޸����{�#����(��c��&�-�e\CQ�D����pG[�*6[mR�'��`G�иq�'��E� !�b>Mn��� &p$,C������x\@H|ʥ ũS�h`G����T����EdB"�վ�㲣HL0�#Q�;�7'�^���p@H$X�=_Vb��&p$*d9�'���S1�#ѠX8ֶm[ $"�����#M㡉��� !��(�D'����bc !�ȿ\PL�Ht�FS( $"�rc $2����#�D�a��Ht�D!�&p X ��k(0`G*�<�P`��B L�!�P ��B L�!�P ��B L�!�P ��B L�!�P ��B L�!�P ��B L�!�P ��B L�!�P ��B L�!�P ��B L�!�P ��B L�!�P ��B L�!�P r��۾�dcVj��=l@E�@��vk $"vKX��c� B>A1\ν�R�i)0?�z��g{ݑ�[e��&a��,���R�@@��;˨��F B>C�Y����g��N�Ԥ=S��^y��%p�63�L�ʺ�:�B����pw�����w�Z���y�fo�������1u#�B"�eq��1H��2p L&O�	���1��$oWX��������_
��`X�" ����8�����a?|h����$Hk�V[D��xF`�uG	,�&�eǙ�KVS���[c $&V�M��|N=@�G42��aх*��I��9���8�׶Rs``��4%��d��x*a����ʮv�B���fj|�������Ź[�/y�b@bN3�~�e��
ï\��!��Bc�}$�%��n��i
��cْ3W/��B��Z�J�e\~��˦�,ѕk�f��(�2� !�Bb����`�v��u�8�����j�B!�ă�,���R�;fbc�a�J���Ժ6H
s@b���!T͂FƂV���,�[)0X(����
	/��	����_�A��#t�Г�Q��Ŋk1�Ď0Se�ȹ�ŋ�k1�@�J�3D��ܑ�q1�Iz�Y�W�z6�B˺�J�>����灕;
�^�a�)9l>)��ܽ���]�F���֪N�cFe�c�.fl��!J��E$9��[���M���B���bm�mb7�϶:����)a� �ƌ{&p?�P �)����c�>���j�ng�o�.� k�VU �O=3Ғ�Ō6�����h��E�1C0���C-�0�Ww�/�3�{��R8t���7i`w��������F���/m��ƍ��������GHn�����X-������e��n��63䘍p�b&3�B�Kw����O�x:�7��ÒGKa�)9��BG��!� 1c� �MW�X�ȵ���J-��1�,�Y_��D�b�J�� �$��J��րf���q�e	��}/�D�������T��;ˋa[�U02��f4���yBW#�Ez�w���a�65�L�W�@��^옡���M
���J� �9��ۺ���p.�����H���%���r&V���#K�s�/ԡ�N�����:zq���`��.�.1fxMQ�+(�G���-��*��@>��!Q�R_���vq���,��CS֩i�F6�6�����h�J��`��p���TD=��PA�
�~CCT'>�rN[*@�km�C��q��(B����K��� �r�B�5��>�1��\k�8cI���V��u��	�T
/F7��O�y���]*`n�r�|B#rnP¹/��_Հ�)f|�U\��x�W�I]�^ⒷZ���,sXT���H5��"��e��n�0;�$Rm�L��W����"@V~.�;�7$��i����F�[���Տ,������`jO#d���bƌ~F��;���NJËQ��J�V����M���	(�]�P��|vUj�0W-�����Κ�e3�d�y�����b��X�<Η�1�j6�2U|r�Z>g�܍W*o��74Ԯy��\5��B쪌`Z�����W΂�=��tW%�ʦ?`��
�h��
Dd���)yW�N�r(0JD3�����s֊�3f��b�����*o��z��0�fB#���X��g�����
>)s��۳`����_���ud��,r�=i�������ʼZ#��vwY釉��e����?�i�6rʐw���㹚��Ӌj����@E�ːf�OZ9ܭȉ�G���r��w'����O��c�#���oҗV=��t.��\>2��Z�N�W�\�`N�ȀI�ˇ�o�~^.�n�u���l6L�4sm��ۜ���2k��ľ[{�"�F˔^����{SJFf�\����,�ʞh�0tk�v��v��c`H$�0T;ዜ��7��c�A.�A1���{7�'�d�+�v�@G�o}�p)t�ʯ`����0|1�^�e|� +%���e`���[J�v�nS����ֹS^f&�pf�`�����.x��K��KV�mSYA�s��t��e[�o�nء�2h��Zz�VJڠng��P6�&������,��>�kP�Bg���ʔ�T��#&�g�#����}�7I�7�?�QW�,�0��w���w.z�:f{���A�H�X4�މd	S>f|&ǌ��e�k��Z����ǲg���+#9��:$�>m�|Z������m���U�&���!k���i���{B�7�Ր�i��Oj��eY+�׿9�Ѷ���ζ���L��%A��M��K�h1Abd=����в��ƣ[���7H�&+e��*�r���c�
�-hQ�Y����j�O��P��#����bF]ƌ���b�+>��!.��0�����-{����ӆ�j��w�5�}�v���U�S�?ۉ+��&)*��)�xad�L��1��r�$���+z)}G{L�J�7�8kF_sh�v� �9w�������/{�^�LI��7UH��yғJ�����f��̇��11rƒd�VA���=��nW��(X�z�tw\�
���:�K"�.3��r�(���]d��$�J-�E�&v�˘��:+�Q\̸�m�-.D������bY����:C��K�1���|��p�C{^#�
�]��͹���W�_�	|ς�ԩ�6q	�?����x���|O�!���5b�:����4)�\�o�s\��'���ȵ��^�y���3��A�����j{�]��n�~��/S�����չ���f���r�/Ǉi����`p0ؔ�Pu|3�;O�?;gT�k�C{J���z��z�����7К2�4��M�r>f������#���T.����V�]1oE���c͌5y3��*��A �͖_�,XXm�['�v��;Ax�ݾRb��f�6ζE˝'p��Թ�_�Gh�E�ڣ��W��I9�O �+������M�S�2�����!�	3|�G�NI������䕘q�Xb]sT��W~Ǔr�'}>f����&Y�
3ȥ��:��Ýޏ��}EV��B��B�m�`
��n��;�����(A f��`e���]m�z���F�¤��dX kr��S�o��!��N2��L}?%޲aH����5�7z���J�wNA(���1���C���qH�sOq�Bǌ�?����?hSǸ~H����1�������$u}�auX]搚�P�?�(���o���ξne��2��ϝ���H<����$Ī9�j�/V�!׽�5�� -1Q�w��o�2��L��5����4��c�,o)����e��v�9�F(P=�}G�{U�<m����y�y���5���_z�bF3��b��ޝ����<����~����˰s�~�V�Э��1B��s�%GwwL�����r>�����*>d��W�
�	�A�|�_1rJ��������ierΘV�o#5� g;��]*��c6[�D�Z�nѥ�Ōþ���mZ���Xk�B.�
3^�>���3�U,9-�Zc��#B���g�\���AgffV������M����@r)ۂ��lƔ�h�j�j��� o��uu�������aS�Y>49����eɶ�:��S������fXr��S&"$6ø��1c��E�"�:���G�b�.f,�b�02��l$���i	�*D9d�fO;�����u+��d�'A zP������ Z���m�mV�ѭ�� g����Q��:�O��7Lzd�fM�z�w�̥8�&K!bG�N�!>f�U����}����˔k��ʝ� T��f�l���$�Gsw�	�{���a #'9W�E��@�)�mGd��/�\�Q��� 	K��s���jv��1����+N�	�T��~�c�W{/jk�ja��iY}���-2W:B�3�,f��v�C�W���i��Z��zZV.f�>4��3�f���Li1rE7�K�M�Z{$�էm@ Q2�������6����j#�&.��V#IXOyRN�}���T
�=�N���$�-�Z��x�E�!�ף� [�k�7��7�p�'9#�܂����VAb�.f��*��q�=:���	$fx4�3Z��֙��\�;Y<��\���l�,��<�r��P�B��v\�2eȸ��*OԪL��3z�M�	�#��J����?Y=s��ڼ>mʈ�f*�K���6zw5��	��I�	6�ʟ���O(��ck���)���=k�'��	�Jz'z~I�Z̐�]�x����2{�]�J�\J��;!b�7{��2�:M�Dsu�+�S�~�:kY�:W�M�ߡ�Z;�L��[:eЏ��V]v�����R��6lЁ:r��kFj%�$U��*���d���k�Z�k�J�3���N�cp�a���u\"k�ui���q�)���z��kʠ��tؓ4�[#[O����ZmgfC�Z�K�cƶӲ�ӏ.�4����{�fumd��.���Kՙ=\��;�F0-��)�X^�t}�P��OM��\����Ȣ�
E�]}0oBZ���+���w��۾֯U���m�J���S=TW�Tˀ:AM��|���&mRZ��ڠuQ2���݆��*��C�?�w��7N�M�������^������.�Ư��}e�@��:/��}�������u��Ώ��:�1C*ʘ�;_6�K��xR�|Z�ؼ����e`cIᒸ3�*�LyF=5�7W���N�C���R�"\&��{C�6R&��?�۟sV�}�-	���'�1V�M�)��^Bԙ�B�C/_�ֈ]�6��UYw�Ab���M�i��)jm��_��a��j��3>"�<=���cC"oy��_����޽c���<o>?z����c������t,��Ƒ�G��t�o��\�.x���I�Gj�b�7Mx����4�txԕ�|N�\i+�:�B\N�-W�Be��ӆo��`ƺjRO��2Z-�,Y�mK�`°x�ZI���O�lǹ3���~����W���G1������\)���U�Q���ڵ ݁f����\��@1JJB�q1r���k,���e�ypT�y��P~�~����>������� ��e�E��Ƒ��.M
�e:���^�����%�=)��1���0�N�w�!D�,(��Q.����,s�V��Hb�hy|]�BG�j��Pw	�F�vvr��2�eCQ��D��'��{��| �
�.T-�[��d��o
��E���}�]�g־_^�ϧ�3R57y�#M&��,�G`G�h�y��7�;f��,%���ޟ�������1PU&FҬ^O��[�H(�Rh���=$7��2���p���d�s���D�����G[��L&���NQ�����q>U��DOf�|�Ơ#� b�:������dm�����m,�j��
�I����nd�u�y8lvuW�?v�Ƴ��\��\,C�\!�;�`J�����QQ���i���8fH�ɐ-�gۂ��QIE����HDi}�j����v�U�&��e��j>;����d)@O��
��S��I!������r���\^��42�cƕrI��� %
j���023|�$�!�f���:��{��*�8��}�\�K�@�Y�u��!��
+囶~U�����S ���{� 1C��/��RO��)�^�"�>�r��x 8+�@A�T:D��I�.�� �f�v9�j�Ev�ոo�`,�����"+#-�ޭGe��y
!O	3T@�����VEƃ_���[�
aΥ�J�Ȩ(.�k��\a��bN��B���e&�燐��~F{#���6ގT
18Zʲ�',�;�BH�T`�ZOh��Kn�����*�A%��"�KM��RS��O�������e�r�`���Q.a=���W�
��	ʭ�"�������vr�ZRH)�c�1Vh��H:�v�W�&�l'60���Ul�`�g�̧Snߗ!_2X<�z D����3 � &��ځ�!IzJ�V� G(��:F���˸3i�{+�"Hz�����_��C�圽���	����@�L�5t�Hɑ�oR���f,k���Ѓ9 Ro/MM�	*���8uU܇V�����?�D*�vmSyn����8j?V:9%	tZ�^�"1#%ʓ���>f���y�X}�g1�;�֔����B{��ɘ� ��)�(W""t��)O������żK���[��+rh�� y����m�o��:4No?^H{���wQ����N��Hl�ǌLG5��X/��,1>�"N�	�L��e�⡅q�@���"N��B�!��!��t��([C_��#������]t�C�.��d�L�߱��������B�1�S�ƌwV��tlh����7��1��������|oIO��Ȕ�q��q���$h�O=�G����3^[���"\�(��{�qMWh�Vab���.*��k�r��������3Β��ejp�J@$�|��+���2��q�7)B�>fH=�;C����y��G�.��X��3���2��}��oF�0����S2�x� V�4�B��	"�"A�2J��`�ͧ�L�ʶ�ʹ�a�::F�c'1��Dr�dy���y������^ه��BGϾ�����3j6`�Ck����N�޴��e��!�?ه0���1cP����e)'=��l�ʦ�65w���&�Z���0ϗJ��޳u~�4i�L?�&�f>�S~��M\�fօr��3�R�q�5��CQQ�-��.{��+��y����ר>4l�q���t��98}�\��9�5-��s����/4,Z�H�vZ�7�x���1#��c�bFZS�"� 1�l����V���^d����+aRw�	J�`]K�=�i�������/����%9�f��۽J�C���߰<���c����/��v���޳	|߾��e�o\Z��F��#��_	�|'P���ǌD.ftk,��ŌF��K��=���0���׻U0�[?1��z��b+����l��̞���  { �p�[#[��i�݇��9��^L�.L��g�1Z�p1��/cF��۩��6���<���^K9W����7�R^�&�d�ɤ�K�f�����������3&�@�2��-��r�D�~:���͂��Ō��\�Ō���u*9Խ���y"nX�Ōܫ3j�fl���P���?�֠����^�d���c��Kff�t�۸t}�h�`�O�&��[�;�%Bb��U͝�����m�4�eevʀ)Co/���IǾ�6
3��J���	��iXsL�
S'����A̖��ɋ��G�y�\�n-�}��l�d�MZ#_�3i��Bb�j.f0f�D;�1z��(.f�qJ5F����zw�vaZ�e�^���}D�36z?=M�Y}������b�1mL#�^NL�ZO��e��i�$rr�*ʜ�n�8��If�/8�%V'���7BV}�3�׳���K�Eq�OcF����n���G:�3�b��&p�k�Uô^F��neWq�Ig��_k�M���Bz���Z�4��^�P�ڹ~p���i�ܢ��"��-��lN�9�T����65�y��1�I�C�$�4���4�&�~���3a��1c�ʔA����׳u�l�Z̘�U��e�	\ �`�j��0��x��0��5����u6���4\,,��5Z��F�X�P&eÕ26T-c���l����QZ��#Y�m�oj���0@ș��p��i���у�=9�8V �/2Rgʭ�	���.fPl���Z9��ar1�N����Y5��Z�y� HsУ����E ��'�c�܍�%����,����b=/;����x��
`�:���ë�2R��=$7�ǌ�"���@v��0u�f���hј����j�$z����l�n�ۧ;$&ā�����z�`�{��/�������p_C�'��T�������P�=��#�W���
�ޥP�aؐ�п�� F�v���a��)w���>�)Θ�0���k�(�?U��|�C�����Qb%�P��� t���e�[�� ��l�zX�1Хs{���"1��A�������O.�C��.0rm+��`��L14����>s�~��
���a���SO>}��E��a��� v��e��'_��{�I҉�O��-`�C��n� 3{3�	��3Pa���$���bH
�N/S8Z@Ã_��$��8�W�.L�0rN��?,����f���C�@��{���0j�h�$	M)3]��q,@cF��GHn�����X��e�XY
�V�h3C���-f`!0��!ˍ��I�S
�;�c�wR��c�~���7_���������W
 ���P1lt��(*pky��ѕ�+����.���ޠ��*fP���*HT�!F��0ZrJ*�!@�����R����J�D��I��w��+�����6�Y^�ʮ���YjQ��}K-�g^
Tk��a�wG	�:���mSaۯ;a鏫�����|7�j50p@�ׯ�軣1�Č�����2x )p;��|�Z�0Z#fh�4tӅB'm0��"��)ᶩu��e0 8z��amIl.+���-���1=L�Y�ߤq�������ۛ40s��_�n"�J�W���K�v���_`��^�n�~M���faVݺ�YN�5�z �껯W3�i�d� ˃��IY3hWP8�� ��ZvMT��|ЃC���:�(8W����j�vF�>\
�Z����+����A��i�ͦ(

�� ݻw�����w�	���'7�4ܫrO��<2Mn׮aİ�|ŻY ƌ�.f,����E[��E8W�~*��W�I`@&�r��:	��p�Rb�%W�����Fx��I�g�$w}�_	����Պ�;#����x��1����������#��{��	8y�4$$4�{��\8~\�΂-SS`��!P/�.�K0fxI���V��t'4R)��>�?��i����j-w�+`~��Ċg��_�e��J�==SR��10i���G῟/�«E�ǲ,���a��qso$���/����힊����>)Ɂ׳\(�c���6c�'�����Ւ�_L���2�e@��(�T�/ظ/|��Rav0PI��p�B#��m)���E6���\(w���
����P�?�
o�5B�z����fmS�k��p���7o
�3�|k\�����b�6m&t�։/W�t�:ciY�UW��U1�d6�-����v�;�FGG����.|A�����k1#��ѯ�[5f�4��ȭ�me�((���8�)��R*�E�
���#J���l�bq0�t֔/��'���7F��8��J�q�|�yV�ᔩ⓫��9�n�Ry[ߌ���v�k�q�*���i<�^����mʕæ���+�϶��M������0�)XyD����m�㚕��Zx�����=.�f�æͿ�@5��/|���x|&o'����z�s1�C�a�Xu��*ak�ƌ��c@/���������<�Xf|C�[�����'2L���H�~.V���xk2|:�X~���+�^�����G��7��u/�#c�ȭ�āS{�C��Ke^��[X�����Dy�ˋ��i/���4r9eȻmu��\����E�R�Ap�B��W6��q7=�����0C�vA��dƧge���~:��'�@Uk�<��}��p�,R#���{�������\=+Y����:7�N�Xr@?Rt�h��)��)�M.�Jg-z'{��}�W0'dd����C�S?/�x���ac6
�m��6��mNOE~yw�t�ľ[z�"�F˔^�\ν�?%#�g�\��keeO4M���^�RO˜������*'|I��t���X�	��
����?��'��"3}�K����$�qVhc��0;Y�׭�,dؙb)�(���2�zZ���2~5Dƍ�u�1��VdDx@O��K�y�A��{�٠ml�b��~�X¯׽'�����s-bFBD,tl�Z�&@tP��j��^8	��o�q���2Ѻ�Lj��`(5�ßg��6@qE��8�	ZG��^b�;v��fO_�Ν���I*��/�&�m�^��Re���b�TV�}ǜ�;�mwٖ�ۻv('�[G��JiA�Iv���e�j��oX1{���)�c��.tvm��L	MU8b�3ඈI��c�C��wl���I{�ߴ&.���a�s�,��Pd���;�jX����t

ʸCZ\AAn1��� z4}�v��)��ņ�Ҽ]���r���X��7cFjl"����m��{ f~�������[q6�N#X�ܻ�Y���t�o�
F~>��쭲��"Z�p��\��[^�X�L��we$��S�Dާ�O|�ip���ƫ�\%o��ȴq��aS�U���o��!��������˲V|�sأm5���moϝ�9K�u����]P^���~;y �K�Wk����=������j��+j����|�Ȝ䀳�"�����q�j>�rl�y��^�kߍ���I�Ԣ��yJL����*�!���/̓X.F�?��?��y'o����+��m���V�A�r��
�*.�Pۿu����ӆ�j��w�5�}�v���U�Sm��DA�3IʊQQ2�`d�L��1��r�$���+z)}GSz�J�7��ތ~����n|��:0�n�uk�_���'�����������f�B��;/Mr���N샯v��EO���/�	Y뾩����#��Mbq����C1����ga�����@����5�����k	W1&��ΐ���mx(�1=��О�H��T�/�������ۯ��g�[��a���p�Rq<{Fv����m��?U���m��o.ɷ�:.|����ʿ�|�'p-�6���f� A!��ſر�O�d�qM����wpjw���߲o&��<��}�'���n|m�YY$�\;k�ػb�
�o�Mkf��k��PWyl8o���g��j�	�uq���~��	�����e ���4{�q�-Z~g�����7��ߘ큻��;�m�����(e׮ϓV��jF�G����.�r����	�K�}���;���յo��j�Rh�-L��-�ug?��Th0�Q�U<�������j[���	�C����_�w���#��Bo��šK�@�7�gD��{8׵u2
Az}������yR'�6��t� ��TV��e�)e�S�r��8�v�/���V��b�JCʌ'X�D�q������X!G]m���2d���/�7���8��s�����T��n�b9w#1��VRZ���;�?�^�Ù��!�!�CZv�:�p>ƾ�t^��%�9�� �FCRd}��4��s�a}n?g���Ӫu}M�����XX��;�;�;����32F�a��K����,���!��OKi��0���C�M�h1�?�����ᕥ��z��SIq)���q�TC.\���R~B*7�e�X,u��$1z��`����>߾^�q����Q��c���3\9s~Y����^�����Z��٫��Un��6zAV.�Y�>���g�yF�`�a��0���Q��R�w�I��Xi+Wی��b~�;@^�����o��{8�B�Zϝ�F�X��q�c��_L��R�Aj�$P�|��iAq1��b%K���+$#� c�<���!�k&���=���|��}��Y���~>�������tZ��|���	�>{�U]i��q!<�������X�I����ޤg��]��NǤ�\���i׃�e`k%pٵ��12��J�Ŷ�Ý���V���O�@���ݽ/DYA��QW�.���5�����#���/�0�����-�[��b=���kM�p�\o��`����;����/s��w���gRK�l�0�mX��,h���[�L=��[���L�ݤ���-��.d���C��*: I����w �`�|D��9W�E��@�)�mGd��/�\�QW�����>g�Ȫfm&���ֽ�����;J���~�B!�(�����Y0�UO�F޿YgX�ok��Y~`4���]�@������ʮB��m���հcµۧ
/:}}���7�;�)-F��Frɵ�Qk�����$J&'韮n�j����4Rjk�
��e
��c��S���c:�>��'��|�ʃ)��'2���7V|l^!���`��gM#S�&F�w\(�o����I��L�J�y���ג\�k6Bc'��Ց+U���ŝ&L ���BU
���q97lȔ!㲳��\
������(u�@`�U��N��ꙫw���iSF$7S�_r�}��걅d��s�����"k�׀B��H�q2�Qn����*������岢*'��e,u�����Wʧ�|uֲZu�N�ܿC�v4��J3�tʠ7g�r9$�eOx�_P+��@�B��_�Z���o�NMo�b��-KC�cMV�vӴөu;�1��tҷi�~�Z�~{�����/!��0dRl��F��˯PF��{�ֿ�^H�=����_���w�����h.�ܙ6�i�L����z���˅�-}jz��
�fo�F-W(R��y���^�t�5�	���R���P��܉�2�Z�	j���3�o 7�MJ��R�.J�p�'xCi����������d{��g�!�؜�{���B!�}�����e���N��٫� H��y�~G/�|��/{�V8p�D��}�x�9�v�=ʏ���^�$y������7U���e`#��!.Ɗ�S��2}�����\�r�;琩���T�������D���I%�����Uo�~K�?��u*Lsi�0��K�:!S(z���#��+�f�*��7H�2�I4-�<E��\ՠ��63l3\u��,'zc?2������������`��z$�zv�m��� ���h��{�F"��NB��\�7m?�m��}Vs�}�W�n�7�Yx�ÃN��q�#>{í�3[���I�rj�h�R*�o��6|�%3�U�z�����j�g�*m[������
�>��4${ǙS��]|�̍m�+YOΣ�SQl�UW�P�/�(
R�A�Z��@��GE[��a�X�%%����J_�p���e�ypT�y��峰���n��#���:���`��`u�Ow,�ٕy�b�D��!$//y��	���F�u��>��_��}�(,��K���h6hޅ���PJ���ዧ��]��,��<�v>G\��u����� �eA�r����n?ef���DF��$�#c�}�T��	�6H?�L��|�ղ���:���	�e߾�ۑ$V��ł�%�c˚��,�M�y�h�z���O�o���M��ބ�ʜ/kp��Ln���C�`A֙A!��-���jX����.XM�]a<U%aRa$���@&s9a��)�Rh���=@~�%�.�}_x�,~w�_Kq��o I~��w���#ӡ�B�j��%\M��Qa1 �o��c�����.8�M�p�YY�ԭ�L�
�X�F�=!������v�U�&��e��j>;ĳj�PH����0��X�!�0@!�C&��υ�u��Z�(�8������
��Zm- �Y߁�]&WJB��*�[��+g!I���#��RN���8I�E6��,\�.�\���~�ոo'��FG�U{�[�G��B��!K�!���QQ\B�B]����2Q'tz�m���L��O]Ϳ��0�he,_���sG��B�3�����*�A%��"�KM��RS��O����u]��+���)#��-����T�A/U��i:B!ቦ"���^i�X `;���"dQ�f�Y�ya��ܙ8E��z69�Bw/L�"�J�>j�-|S� v���1�χӑ�`H:?tL!QB�{&p��+��c���J/����A��S!���0����du !�"0�#�B8B��B��*��D6�8B8eAWő�$�$ �L�~�穃����pܶ�8B!���G��O�7�B��0�#�B8B!�0�#�B8B!�0�#�B8B!�0�#�B8B!�0�{ItP�UZ0��p���Ve)5PG�־���(�~�3J��\���A��%& �Ii��?>_|l��}�q�����}kB*�@��)�\�������
����Sp��b��'���~gȱL�B�&p/�1�yx��@Xq�W���Z�1�UO�b�4��}����ŎUN��U���O._{�X
{���������e��G3�3G��Kg\��d�A���!� ����x�mo�=���'
�;[t	���>�}��2�>�8�z�(��ɉ��6�;k���
<�Cȟ0� ;��g�V��C�[e�rJL��c9W+�jiM�@����ۿӞ��~��o_	(p<}_:,xt
��$���[���K�S����.�-c��*�$�=���Y%S@��PW���w����b�B~�	< �����ݱ��E��o'���R&�S:Û���V��࿣� �Bl^H��
��2�x�_�����O�*�(
:�5�pm�[e}�tG#Z���O�������U !����mV��������֢+��OXwd'�t��u�k�״�	��sG�&X���=�=��%{6�p.��h}?ܗ�
!���n��m���ކ3ӳ��L�{?
c��H�B4:���0|�5o�Xr�S&I�!���nA�i�f���~)� �߅�+�=�Nj�?����EK��#�5�x����L����:�;!X��4���c˯�08��>'.�Ծ}�_0�yXy�7����Z�ۑNkq�17V˕|��H�M�F���@�=Br[Ww��:H6�^�m��p7 ����~S�>ʗ��M�B�+�r�q�V�	\��5������BlH$<���F�q������~>��ofwG�F�\=$#�\� ��� �>�B��﯄�ݾ�D��I��T\��nAtu��G�l���5r �;p�4�|��<�Zt�n	-AN��1�d���;��LvkB�ۇ��V�:A�Y��Z��~7�-&@H�H.�?�q� ��	lB dY������#3�݀�u�L��e)#Mޤ��\�~�Mo�1"���!u�h�V�Z�l�Y��Ǜ��1A*���* ��8�C���=�2�L*��M�*���}��g�|��Ua5��S�Y��g���1~Ҟ!-���ݿԪܜ+����3��7)��S\s�w �|8������y']ί�j���XW{��}�ulB��r"0u���l����A�ɵN�đ����d R����`G�hS�	�o֙�I�G�*0��C�H��[�7��,8/��'- 狮@p��Rx�$n9}-t�k�!��/��aPa:
"�@��痍e��n�0;�$Rm�L��SwO�41k?=;�_��4���G@� ��M�v��<ھ�g�R���H�GR��#�U6�`�����vC�.����==1x �#��6����J&F�[�&�QN��R�.�V�e���Uj�0�f���QHgM��y�߼~�pc�k��cl�T����g5N�*>�j-��q��+�����j׼�@�W_�ro"gQ�r�

u����"!sPWUA�y�վ2�f�Zw��pM04�������}��+�{�>��Vy�}s6.���ݡ}�d���x��=��^�d��O���7 �,޳ѭr�&���G��ٲ�{�/p����-b�Q�r�q�Ӿ-Ֆ)��7��+�:c>��?��N\9��	�M�Y+JΘ��e��7dn������>�a
̈́FJ�s�r���[��'*�s|r9����q�J��ل���ud�P���8pj/}��z�̫U_�`w��~�(�~yQ8�s�$kjN9eȻmu��\�ܿ�@5�/�#\������Z��ݪ,�Ҫ� Hm��Es�}?kƽ�r�%�%E_Z<�\�$�?N����/J&D�G���P-�����8�E�w����p�de�C��72�ˍ��!Q7kޤ����,�+)��<2�y�\�'d�Ӵ��Wۛ�@arp��T:k�;�S\�s��9!#&m/2��:�y���,�8l�fC��M3�fݾ��5�_�]=�2������2�g�\(�������3W.u�5���'�&��A�]��eR�K�W�Ju�
ҥ�r�� ��œ1�
��x�t�"�m��z�����Ĩ�>�On��h��G=<���Y�C�h3C��'�m^�֓������6Rs&���X�5?���������;B���k�$��@�w_{x'���?^�*���ٱB�����oֺI�����C��蛏)� 'R��c�`5A!�Y�{C����m*�=}�:w���$��L�Ӷt�/�z��{�j�m*+�c���ζ����ۻv�&>8��>b�N*����ʾ
�?k��oX1{��������\ē����c��e���7O����0d�c������G��ͳ�ݬY
L'����>x6�=���+�ɤ4_��(�PRQ��j7s ���������\n��X�����~��Ď\��0v6��d2��Q�y\f�.�a⋯��{LY�_@w?��j�����,��we|���C�!-p_-����7Qe/���:u��]ua���T���hz���}�O3�����m5��� es�kT��w�ݍ��V-���ھ>{抏¦��V�E����X��ڬUUv��vى��g����d
��ؙ"�c����I�%:�W�RZ�M�!�ĉ4��lc<-'�1=��О�H��u�f6�FV;�f�	|ς�ԩ�6q	\���s������"���5b�:� �B5t�Z�wżw�Y3cM^Ì�r�U��B����=V{�Э�\���ܝ 	��a_)�Y�z���B�X����PeZm�@S@ �6�����V�6�@�]�� 3k�B�Z�:���edR2�S�]��4�n%�/&�4��x�UJ$���)�I�UrB�Z��Cs�*��ʎ� ,,�Ν��[�P���32F�a�f��#��;�Y��J	!�PMɭV2a�!ʢY���\��3��,X �5�fS�>� �\ʶ��6	R+m!�P-���J�k��c�ߕ��m��;��׭L+���A1��{_����G!��� )=������B(�pH+#9W�.���@�)�mGd��/�\��D�Ndd���U�B!T1rE7�K�M�Z{$�գ��z_��b0w7����M�C&���H�	����2��H���V�6�.*�
�=ᗓ{@-�6�P�f��8�	UT0�=~���ߗ� 
,du���]���������L��f��O��Ց+U����|�'�(�g�2�`�p97l��_\6c�����2�w}�:)J�,Xs���~�z��]�y}ڔ�)j������~���Xq�^�P`"�𾼪RlӁ���l�+
��A��O���e��\�6��fJ�h��W�R;�dʠ���V���eOx�_P+��@�B.��JhI�F�U:5�Ɋ�+�[n�:�k�J�3��)TBy&���͔�?,��I��\��ҧ��k��m��jd�r�"Ů>�7!-���g�8M����o�I���P��܉�2�Z�	j���3�op�5i�Һ�����a�9B!a�S��2}�����\�r�;�2uP��ʠ�2��������2��|��A��������oI�}f�m��h�/��IiA�u&B�P����G�5bW��<vU֝o�8eh�hZ�y�Z�YN�w	Q_�V(��BA�`��f��f#�y}f�
T�r�*T&�1m��Kf��&����-���ϒUڶ��Q�B������&��q���g8sc��'�S�HT�[���/�(
R�A�Z��@��GE[��a�X�%%����J/��鄸I�ϩkp�Q�;'�!������K��P���B�}��H�eX8���b����e.P�JIL-��+W��Xm_"��BB���=�(1�`��u�p�N�P� ����P�bAՒ��%����*x�^�1�r2O^�������H�4�$�v@!T3��H���)�L&�	ÔR)4	��� ?�5�O#.)�\?	������:x�a
�9{��<n�BH�0��X�L�bk��o���Yg����l�4B!��.bG��;��V�R�Ձ� нu��\���c�&`�&N}D4�ږ|���f�[!BH40��T}.���y>^��(�Tt	����ִ3�U������V�B=Uj�,�6��?Vj1�#�&p��!p�K$����K
!��݃^x���2���SW�~��Y��%k��C'E����'m*+�_E�&�vG����'X`h�:`��e������eJJ��E@B�^ccY�v�4�����؄.Jdv�D�~�4�3#�Ii�8�nDS�e'4�s�$;W�q0���Fv��������^KN���љ�$���o]��Z*@�v��f��x�ߛ��o�n�|	�Hڬdf:A���\B��	\���
�������������ٙ�ْ���&bÊ��g/w�z�wV���T�z'�x����G�)",����2�yV��n��Β���׼6�<;;I�|��?��	  �x��PQL�&�E<��5�o�B�4g����Q�ղADyz� �u�堍�%t�%1��,/9I6���3�����>/<J�����q�i��'  �x��z�c{�o�])Nݰ_U��Eo�K����Ϧ����u�K3H#�[�IpШ���r��g ��@�Ǹ#N;�<�+��u�����`��+8Ь������l`��  � ERmzơ_h�9��JH�2V�(�o��F�+9A?Uc� @s� W����8p$i��)f�|Rp�{�t�YMUX� ��@�+P��8  ��B�  (  @��   
�   P 8  �!�    �@p   B�  (  @��   
�   P 8  ��Y\�7X��Z�QSs�~r��T�u�q���:mt���{   7NE�Vc��:#eh���kH�q�QqM}kċ4����Ǜj��8���P�h�5� �o_�{=�Cu��,�j��   "eR�t�9�.��'�:f�u$��D��i0V^��)t�9��U�7���Q# ���U*�Zʓk��1Q�n(Ex�Ѩ�T�g4�{EG���&  �p��79��ht�T���==�֑�Yx���  P���Pj&ũ���Q�F����֎^=y����  J�T�~8�-�95)�/nTb���T����;r��T�uU;��j6�\�V�%�8����Sq�`J;�Y���|^  ��,ո���.��rH,�>_5�H%�P\���k��2��W�r�rz}E��)���'�s�У��H���@[A�$��y���.G�!���R����g��.�6��e{����H[�>!�5,�/����ǩ�  P۝RF��i6?�r�q�^��^[��q��gO�w��`�����7�y¦O�U��q����ݞ7)??PS=��l��\�f�9җs�x�IWY���~�`�p6U������*��0��L��@�y�A��t�Ko
l�f�$  ���7�<o���M���>>/;T��+�S�q���3?R_q�J�n��%��{�k��Q仗���~�UW�%~���	U>�Cu���3�,�5�Mϛ�4���&�R�Zz�#����V�_   ��(����<_��x���y3�������o��7~?Ԕ���Q����_W^�����ٖ���e���G^�Z�Ҥd���E�X]�@C»ƂYVpSG�~�1�36���tAK=�q􋣊   zL�*eC0.Q�yW�ߚ7+��`����Ա]g�'/s߸T�7��]�~N��f���z�o��~�)�^9ol��r՗3����ϟ���o�}��22��!qV8�¼�C%��m�L�xR�B7}�O[������y~���kH�%���Ey��6��_L�{�2���Y.%m�U�k�����*S�4��E�t��nK��$���/��Dz��J�ZO���N�Mh2A3:�r�س� ��z��������O��wF��~��R�3�Ԕ~��t�����\��y�\O�㿖|�7v��صx��"������=���/�}��gM�� h��]�ic�]�-˞�<�Q�y3�N�gg��7w's9W�N�z7�k!�2��_҃,^���'���]�H���K� � Z�T!��\e��c�ާ��e�6U�k���̭WX��mZ��Q�0���$����u�ΙՊ_d�^�_}+]�m0�}ɻ��Я  g��CO�r9�!3����w��aY��e�6��a�ܜ9��̸Gԩ"���Uq�H&nm��P�
�Y�����B��J���K �s	ud�ې�G����n9���"��pʆ���Y-��e*��|��.9�%�+ۑ>�N2�O  вյ���n-=��|ɋ�L9�ò�����Ν��=ù�6�{�p�<S��R�Qz�F�k�����U��&: @KWW�e�,�Q����AU�Z��v�P_ٰܪ�#�Xx�&�m�ֈ�ͭ������  �\���n�>��}�j�8��ٯ���)�(�I�~`Vv�&7'��u���y�%�α�ގ{  -�q�3�	B�^�6ݥ,Krr(�>�a�w���$�T�v��PoŹ� 7i�c�t�x�I"����җwGr�=�1�^��� �����  -��R&tӟ��K��կq�y�(�Z���V�����mߐvZC��)c�rF��u��3���2"���<�d��h�c���7c��Ƽ���7��3?��F[9@l�yI�B�*�8r�3#Fp�W�'�76�R��Ǒ���yܝ:(�	���e�<2�������1�=u�ER��J2�7�X�}���9_�U&d��x���&n��	%�,�F�S\O��[�Ԭ����l�k�N��]gXl	U��祭�
R�Q}.��I���n�m	@i,E�@�.�F
p���z�C�Ǖ1P�i��X7�uM��[l�4&�K� �Xy^�Ǭ_�M���♟5h���f���|m��ndiR���w��N��Xt���~�W�D�������5:���vqO�����_��Q��]��`�*��t�,�(
4�(������.& �p�VNx3:��2qӁ~�&�ݢ�VVӸ����[k�&�sROy݂�K�ù渉�o��}�$h���6�EoL���ڿ]y��W��R��Y>�;;���/u����|�҉�Fse��4��	[Oyl\0k��`�X�y����Co"�1�V������dE	*9�5�n@��{DE�w��O�'}T��t+d��*��&k`m�`R��rsʪ�g�֟�8��x���ʍ�4rpkA�nw��/����:�)%�ͦΓ�,�������y�9��Y��-��2*�o�_�&��a"(��c4�EӦ���j+�x��D�)"�_�V�%�5Zi�&U=�(���E�ȯ����� ���O*e��;-��i�'���x2�#�������d��+�֪2���'�$9�J��(���Qu�X��Bk��f�C�۝��x�{|�|WR=H����e�~ �4zc+�i�k���H��ؼ �1�W��M�ީɱV��HYqoJk��R�αf�֤�+��/�-���+��(~�V�������#�  ��-�
��趤������#�� ��y��ҧ���j  ���������Z��iR*���V����T�.��@�L3�fJ�1�.�V��z˖TW����v���ތ�j��BZ���N��~>q���\G~˘��R�ꨦ��hBb+�k0�)*�E�;��T�}ΰv[�0	j5-��tM��q�OidAWXXH$���=�^Om۶%��ؠ�Uڪ��O_��l^N �|�
���#�Ig�k�JKw��T
jV�� g����8ˣn�j��^lR�}�t���ױ�OKK#A�СC+�Z-u�҅x������&z��lr�ܔ��;��U�a�@m��������k��O�����D��j́��PcC�]-`O�.G�Zu�����?�\���d��ю����������=��_�Nk����[\ݨ�>Sbb"Suul�G���hTx�`L޺�I8@�*���%���F��j�W;�k}����H~�Uk޴]�{�B�gd�+�}�q�9��͏ӕ]��Y�Ц�;�ym�6ta�^�`����G��VkL�J�?��b��:���ց~:y� �ebk��c�w������1_"�b��|RL�l6I�WNj��A��u�� 1)6��B�R��<�v7|�w�:�.�,tٿ�`868�+}��x<�r�4@���v�H����$ )8Ȃlii��г�&�)p��j���,�Y�|UUU�`�^߽$'�? @�� 6�����-�a�An�`�����k�#)))��*++:g����	�5  �"v��):y��=����S��PV[M-�M�6TTT��<X�޽{S�ؔ2 ��a�y�ر��c����Ifs�W7b���Ck.?q�D`Q���r�'�g��8 4K��fN�v��g=�~�t˹���i��k�7k�NOO��<ϛdA޺u�@3��#GNOgC�@s� �_�?3�E�D��vxk4j߾}�ټ)��SYX�&}�/� ��9B�C��o�ݡC���^��F�8p 0�! �Ml��m������]�`qAD��4`G����V_c5o�N�<�{߾}�n�	q���s� �x�4|�PRYV���o�*v�g��Y`��nh���pGJO @,B��tx]���:k����c=�k�~�N�:��!��l��5p �Qp ���
4T �ala�5�����j���ۿ��5!޹s砋�8���g �X� � ��[���b�k�n�j��˱Z:��}��a��)))����;w�g��V�cϱ���l�7 �X� ��X`��PCa+�)yyR6W��g�+�B�մQ� �A�C��ȕ�5��mۖv��ՠ�  b\�&z��{iL�a�nI�rG�ڳ��]��<y��>�<js�懳"lu  �B�7�+�
��v���z?w�ų�]Yx�}�]����siB"�2������?ӆC�F�>Y��k�E�V����� J� obWu���.:'���G=p:��۳�V��c`���]x�w�@�G�9�վSSS�9a�ƱP� =  %B�7��:�<~�i�9�4�@��.��G�ѝ��9�/}�1��̧�3�mߋ��)j��Fh7��Gه�3w/ Pxk���y�<q�s�v�Gf�10l��3��XY!��n	��ʛih��Qp�\�Mc˭���� @,A�7�S<��,%��uι+�<�T�?蒞?�%��6�ܭF��v���%$$ �@��MLP�d�o�Ҿg��ǃ�=J
~&�����ϛ3Vg��`0 (����(���)�ʒDŧ���]ԡw��5��}�Ig<V�E���f35g,������J Px���O�=q�m����~����J5k�����~^���Zu<��rb������"@����Y\�7X��Z�QS�"9��*�z��A{]6:貓��~g��p=z��Q�9��ݽ��&��cҿ��wm����}��tx�q|_T���V���ܱ8  �"�5Rg��Zi���֐��H7�"�������s�'q���i(V���i��f�
��~�������y�9�f�Fz�\z���@��5�]z��׃��cr]֩U8��(�@W�����@��j���$хFk���#��'b�N���nI�+�I���(px��޿�Lێ�?]:�z���Hg���,�K��8�5v�K��5�҇��ll:ki��| -� լY�\#�J9�#�PT��`?����V0+:J�7)��=o���.�_~f�y4�)d-�^�� �2�
Z�/�eh��Ҩ� ��Z��'�:�?
��A^-�����7���5Ѓ�m��)�o���1J!��v��Ƀtč��ZR���+ -Y[���,e���}㏈�����M*U��s��b��U���*IE~=�-I�ƬW���`��R3if��f3�-��'�Xj� �G���ᄷ�����J�*H$Nϩ�ɼ�$��I�0����b����/�gO�X�3��,�f��t��/mym��y��]���.�+B�k�r>9kB����Gx��V�D{�1���sGRkz��!R�a�Ző��	�  ��Τ2�3����^t�c����\��䬾��o3�]�G�����t���ӻ�U�w�,|���U�P.Fܞ�Nr'�'�`��O]��U��MT�%RM[�d�����y�C���8�7O������C��{�㨿�B[m���4�F���.y�~Z� ����Mz�����h�|:wzތPe��|�*�9�e����OD�F^�����,y"�����>��Ȫ���w���a��u�4��E��z}앣�f�-�5����Y��q�/0ƭ�煠�~�5���*I$�O/ �ȱ�aMy����n��]�`��p���̼��G�l�,0���Tv�����U�CW��|K��!���Z�Y����^����I���	�#�����y���5͜��j��[���r��sk�lj ����"  �^z��׵`c���ʲ�5��^�X5q�/�&�'�<�
�G�`��*Tx3uv|3g���)c�5̜�G9ol���/f-z���_8cɗ�i7-� �2:���p  ����z��*o��%{�/g/�gy��;-����UW����%k�*S�4�SB�C'܆;�5�Y����9*n��:���;�}���ܦ��R�5��ъ Т�,��]��x%EwE�E^���[`�xY���N��?�/���7��s��ݴR
�帱C.�ΕsVFz6� �	[�������4A+�\  -W��#}�[��r�ί��=���T�g&��i0� ��s'P�k;���K��9��,�x���%ɤ�������K�u�
�5O�m�ko|�����  p�4!��e�'r�O�ϓ'=���^���)V�w�[W�=C��wzh�����u��+~������V  ���Ŝ*�Z�����ɒm,kh�߆�3FX)7g�G�93�u����9�~��So��V�����,��:y�Q��xh' ���:��+X���>�G��D��Sk�P�
���,�����'������d��Uw }�u��j��ޭX� �������IԵ崺ڞ)=�,������aY�27''��m6�
��v��k�f��q}����\K-u�{;@3c7s$J�R���iZE���C'�l)qY���r\G%��'�s��e���a�E���d���$=�$ǵ,�m�Ν�*g  @8����X��M�<Z��5M���,�����r�O<Ϗ'��x�>�+�Sx�(�I�n���t�98#�ΰ�a|kA{Q�sn���� @sS�N �/R�Ie�2��*���������l����%�����PD}�,�2�I2�#=�[q��G�5e̓����k�LGٻҗwDr�_��zm��N[�� �t����+k�ic�u��Y�&�5RM\��2�c�2.�Dr9��~�bvݳ���Qwݹ���
Z�טW�<�{dz�ߏ�[e���^��?yԣ_�\�J]��|��SG�����$��Fӭc&�|gA=�ą2jڨ��u��C��T����^\�}�q�>u� Z����3�3�\�t�g����A�魷<db���/-�֘k��8����$���,[�u��r�U&�o��/��!�I�Pd�`���6ZVz��g�K�6�#����%ĭ6�|Хu*|�jWN����J  =[l46>-�^�5��i�[�2���K�7�#�ѹ_�yy�-�#!e���׺��_�u��Z~y�2A|����Ȝ�M[��HQ����.4����<rB�ɏ�4fx?}ܢdAri��Ł&   �e�
)�'�=�!��Jد�|�y3�5Kj�Q7�Y>a��%]��D-�qT���ֿ�✅b�
�k���k;��RGA;�ȩ��k� ��/7��<���	�����]Ym̤S4�wz���uL�?�v���R  8S~U	���V����A��ܜ�BʣM����Z�9X��SG_ԊӼ��`�>�`�������w�<���xr�?�^�����{�J)�AG�>�*U2O:�����ܻ7�����n/����S�J%jU�����������z���	�o  8�O���_t��lՁ4!*�����`$�͛z��j+�z��
U���p\j"/�O�����։5��$�`�qhRfQ������?�wVq����t�� l1�-϶�w�1:���o  ������/)��Z�U3�z�t��"pu����/�d��0����_�v{%5G&���^��  "��VI�1�=)��
�	J�^������l�qj..�؇�:�.�ԗ:H��	������ǭGw�ʝh�t
}�  ���VN�>ݝ�&��t�P�o�U��'�_B��b�@i�D��]Oӵ=.z>N��B�_��z�=�����ʏ��M[�4���W��7 �]N�,��>�h!%RT����_U�������mM�ħ��'��å'iů?�O���i'�Z�d����x����c�L���ѽ>�����a|����a��+:J�U��pK2�қ�SP�zL8[����e˖G�a�
���N�Q���͚��|}�廐5k��X΍��/Ϣ����-Gw���F��|p8���<uKns���/}�<����޾ۅԡ�%�<����m�(��Sx��j��B�.:c`�Y���z��?������Q��@ɉK���IZ�z���fv�ª2���i_ѱ:˗;�诟�L��r�Mx��G���[B�(�p���R���5V��\��=~1��s��#�RP�Bb]�k�JG�T��~�~�û�W���"�yW�y�v���Q9_ntu�qR�[����^��s��
��s��� Z�c����t���Xx� �ak��D&��^�1�K$R� ��bp���>�}����ooX���z �#�R�O h^�M,)�J'+K�~���u�SL�,ؼ�'>�o���TWW ��4��
�h1j�2�Q������� ���(>>:b� ��Ď��
L뒒I{
�'��v=O_#Z�{����6��  ����|o���������a��5���с��޹1Z�GeeeԦMR5�Q���Ŗ�` 4�&�����ϗ�D�I{N��+>�7P�fZ�����~�V�q|_����WTT��j�樴K��2!��خ��i���c��z,��ͮ�䨵�Z+K�2��8����5�>�����{,**j���� �
���K}=r�ֹ���}��Z*6RseX���(�Wфw�D��]�����v;�w��h;y�$ (<�&s��ڷ�7Q��?R�֝����5��9eY��n��&-x����� baסCj.\.��@��1d���ǀ̮�]��v�����^T]Nۏ��vo�?��`/��l2��98v����!�cЖ#�G�9z�(u��]�#�Y�@yy9 (΢�h(...�5��>s�Q��hJOOO'�b�>|�s�	kY`�;kZg+��v ��Q�֭)99���YM����E�

�h4��l&%:t��Y;�Y,j׮�Y�Ų�G�	L� �Uph߾}Щb�9�NG{��!�緽�Yv��-PcU�S�N��t���Dm۞;P�}_;v��{� @�B��MiU�<o�]�t9��`�ֵkW�lt�F���k5B�w֬�V� �U���Q�!�����o|���ԩS'R���ؠ5�jP#11������   b�l0�U�v���^��Ν;�lM�5�<x�����j޵��& @,�Ϳ�p^5dZX�g#�w�����s���y7��<N�<7q �C�� ���Ez�^ȅ�^\]Nێ�	,�������XP���ݻwB�M�ڹsg�Ϙ�dS��*���ј� �e�P�v�=4����σ)�*���9_�̤�h�ڳB�/}�`����Y���$�Ś�ق3gNCx@s� �O���7���?�X�m���4j��Z}�9���G��n<�ƽ3�~9q��n��gX���8[��)�B|�Tǚ�k��Fx@s� ��x�u˓�����e��l5�k.��|P��t���鞋n�.���⯯Ӆ�e����Y���'ΰ&l��:555�A�V�;q��Y��5� М!���&�լG_��vQ`����3��|՞-����K��C��[^;~�$jJ�O��T�B��%HY�� g�晳�[l��H�Rg�±y���lA˰��233	 ��B�71�tΚǗ������̰��f5��?B?M�����<����QSb��B:XM���KJJ�3��g�_��]S��σ�cM�l����|�[V�� Ќ!����.
<>��m�q����[B_�E������AM���,���4;sIS�,��#;؀8v����ЍEXs}͆,  �����p�u��u���c��~/�J�<.������Լv�j�؊*մ���v��́ g��"��}��H5��˂�r�����v ����NO�uq�J�R� �A��Xh��E���5���M�Kq�����&j+�J��Q��ҏ�e�]e)U�<��it���Q��p���k�"��}�Gi@�)6�,�>r6�,��VX+��ÿ 4o5OWZ�h��J&u�6L���ܘ��`���K2]nN��E�B:<
߷��VA)����1��aJZ[S�l��H���C���i^��+
������n:YUJ �<	*]+e���!(p̌���A� �W_���%���m��q|]�m0��u1�m[ՠ׎���kDbk�>z}�'���nkT�3����ƽ25�ˁx����(�����M% h�R-�!9�Zi��T��=�ށ�Yx������o�.�/�{�V��vm���vc�K��v��_�G|�-~�~=y(�\j|RX+��fj6"��ɓ�Qⱄ|;p� %$$������}8aD؈���L�~6��T4�k b[G��LiKz.�wR����1���pZ;z]
��
�y�ӓ��N�3(��Н�Ρ�Gv�,ϩ��Գ��?����|Je�*Y��_��d��4�Y
���:�����桭�@NmGZ��Y%2����3/���8je"U�����=�J��W��T~���O��A���9��~��d�̂}��nJ�6*a���»Gz{�8�}�n�f��/?�����5�%T/h׃&���&�^�ͮ���W�d��"{ 47l�ڃ��a����K��J��/��"�W�-ɂ֬�&�,/v:��.g��'�&�?�=��y���g�S+���v�������.G�A�c�����v~���eߥK��%S�?�Ag�93�vgR�y�0)�B6l΃��}�Q���te�A��.�����/7x�@�zw�JЛ�y^��I-B;��ՅG�y~ӱ����Q�+�u����;m��\�Ni�o��|rV�`�C��T�����k����y��v�+w�((zuu�U��L
�';���N�eq�f��G��JS������-n�W��lz޴Pe�s>`?��ؑ5u��F�sF����D�f�b�$�a[���~;�:�Z�{���ݓt��ӠNV�H��M��w���~%��dѯ� Z-�Uz�����X]9%wF��Pe~�`>ώ[���9�`����Q��xܾo*J��7j��Qd�쥯���v����24��L
��z}�+�F-|1�p_�;=o�k�5�,����>ҚJ�앁O,JÚ���aI�`���4�x���>�JJ��  4kQ!eC(�^�gcU�Ջf/�>�k~�|�dǓ�V_h1-2�|T*���N�w�'����7[��ٖ����[��o�fx|�*��d����not�߳�Ņa�w��'�̺ؔ<?X_��S���$�������d  �^z3%���N�_�l/�Z4{q��]c��&���%��yr�#��y�M�eW�
o��΀��|�}Ҕ1s/7'�I��a��z��6���g.Y��؅C�	c������   y\z=���/�X�����b֢�-�n�c@��
������x�:���u�o��v�vW+A��㦪�^�Q{�m�^��3�U��X��9�Cw�1�d�W�"m  !��y�}�e^��^V|O��Q������)�S��M;�v9���G�+Wo��N �=�\+� �Q�;���r�ʈW�X��qe�3Y��aH�slr~���lD Т�k��1m�˾��̧�X<�S������A�|S	�q�c9���ʅ5���zOz�%�K��/I&e���aH�si� �±�\(�~�Gr�O��3_z�%�K���S.� ��|��������6�L��Ιye/�  �3�1��!�ΐ������ڎ)���+�����6g�=�N��.�J�K2�j-!WOШ�  -�PǪk��=r���S˒m.�/��xnX{3����Y-'�y���Vz�処�Uw }�u�OJd���i;�y�q	�}�]b+*�U��k���G^��$  -���-����v���r���y��q��,ssrr���+���C�	��ac��WzX)˵��P�}�	6�FG/���9�2�T��������66�i�����v#����7��  !Tױ?�N�L΋|_9�������@�rM����Z�>�I�Z�E�-�1���=ԹS
�#�û�N��_~��,��l�z�z��@x;=n�rt7U�Q�V��]�e M��.zf�\ �s֑f��Cz�@��I���H&VR�̕'�S�(�I�F;�mP���6,{�Z��(�9��wl�Oʅ�{�_�V����))�BS���nx5�L�@�Rh_��}t�����&]{'����ұ��%�"�B�  �阔l��`+����.��&.'�"�:2{�����G2I�hG�S�� Ϛ2zb�Vo!��5�3�el�������7R�ڠ��:mu�{Ē�/<�{�Rz��sN?���m�''�dv���>+���V~����E;����
܅  �X�sV6��-U����ǾF��p$�����ٶ�f;���:��/�/�����7�����ԛ�#��6��o��Qs�p���L1��!��P�7��I):%�<�ߺ���:�;���m�Ц�;�y�����@�gX��  !l�Up������'F����s�1�G륷L ��ԙfز��lYβc�ʄ����dښ,he߈�m�/μ���>K_\ڠ�����n�Sk�7�X����m
�NԨ�OT�s�=��5�s����kheY� �Y�*�����s��Nb=M�54ut����3iL�>ƸeF��[��J���g�^��%���cM��C~�e���Z����5]\hI�E�|�-f.��kF?9�zC^������@�R�t����}��H������ ��2aEEݔ��|��u�۫�4fԂYV�sͱ�Fe�3}jkk9t�4�m��O]w�����}��7���[zf�����(oR�$��Js���d�r��x`��%AGݍ�tÐt!�=q��:��u9iuu	  �)������S�&x�e���^a��>�������YK��:j��2�:�G=�F)��Vg0&k��:M��ǣ'���������y�<�T�o�w��K:�뗩�@�e0���ս���Q��v����Nť�B�t^g�o�����b2  8��Dz��=�ށ��v�2���>��z�~��f+�-��oIy��$hڦ
Z=�g�B}�%���&���'gWy�?y}��|g�:��䒦�饣��e�������/攂4�65���;�}L  �'͓*z��dR]�gVaL����6'�e�9��NK��e`��ݟ/l�����i�]9�  �i�d����;�2-�J�� ��yi^����o�zz�\z���Ft�m�d� ��cS�Y~ܓܚLj�Ơb���,=IUu�s�ێɶ  �i���f��	i4�h%%RT��A?۫hyEr���  @P���}WYB�Z����D�cd�\b:�ٚ��x��i�Rx+��  ��U�)<hN�#�xg��2=%
i��O����Z@��Q��@ɉK��9E�� �y�*�k��G6�M�:��ϥvx��*�~B$?蝹ʗ]�{�~��  -l�K����z�{F�H��Al   -  B�w�G�Zu����\� �~	�dX�>Է?�/~ZM����  �а}���WG���lXB^w���!�ׄ]~��_�B�  (  "v|�A����a�����A� @�
��p��D8  �!�    �@p ���*i����{�(,+�h0ӵ]�Y�`�	��ȯ�	 ��?젯6~��s�Yd�fk
�\sw�e����   
�  h�*����Rg�QA��  -���h��5u�L	�  �@p   B�  (  @��   
�   P 8  �!�    �~iz��?�]���yD'"�  ����ԦM�˫�*�� � Z�r��z����2O"�]|W+��!��q�>�z=T�q����;���Ƹp��ɭ���O�Y�}[)�� ��%���ѵ�2��Ⱟ���/齍K�._d���R�*u����H�%85�^�!^��̧8�T���M��b���"S��~d��V���������������ѨJ7%�Y&^o"  �B�d�C��j��0'ѐ8+��1�0�#��'b�N�a?ث��0)X��(����Q# h���'聼W�,s����3A�q_gI��-Iī��'�� ��~��[S���L�*<J�<.y%I��,�[g��L �L���;-�R�Z�/%3�T����������#�O�M7���>�z<κ�� �4�tFz@
o}��o7���a��?���7N�.;  ��N�����Ъ8R:��(nT��bV�2L�j�@w�|b��]a�y�I�j.>Q���uO�H����OS3�S��C   ���j��+�mR{�����DQeT��I�ƬW7��b��[�t���E����.<���ݮ;�T��o�mw���=r�K��/:�Kr��U��}�.�W�`&o��AgHu6���zS��  ���Q�3�5���l��Y}��9K�ռ����>�������k[��	�&�@�	�>������'�^^���}�E��d��Ɲ������Z�;���r�)��DA���-ntT>���y١���|�:b�P�W����88�<���A?>u���@��6���B  h:�V���I����d���;}�K���^��Ɏ[��}~��2%�5�b���uu�_W�^�V�sA���_�ߛ�ǮZ{�5m}�F�I�>�oCU�f-X�krg���L�v�)��^#+3B[����2  ������|����\]~��Kք{�Ϧ�MsM�q���%f��Je����ʷ�Y;{��`�C�y���7[�O���jkb�E-��	�-�isu��	����.�K��q�9��*h���D?٫  ���L�|����VW�oHx�ț�x7i�}�Z�-�<�������(�"Tx3uZ��ť��&�}g�%�9ol��r�3|���/��x�e����c�����  ���֐��+��?{���^��Y>�<�u�@��J��f[�?��������;�\����ݷ��J��丩j��_dw��u�e�w��eV^8�{�7�LЌ в������˼n�����H�㨽�����'�Ԃ,s�
�N���¿�W�� ϝ@���:WH>J�;�����%ᯐ��ί�&k��Cj�cs��w׳	  4k�4:҅�6v���Ĳ$��X9gea�g&��ez���ZƲ��ra��.���I�x���%ɤL�~"=	v.��"�#�E�ֳY��S�:@ �̥
��a��}��ʭ���/=���{��/pG��k�g�}�/��d��xB��ye/���J|>��{�,�t׏ D]��E]�F���[J��� s��9DO�}����7�q��S�o�)V�ϙ�mΌ{D���8�9���d��Zv�:�Q!���H�؆n�uԮ��k��g�XuM_^�G��qsjY��%��W�u�S6� ����h9y�ȫT��҃,?4���郏��~��sz<���x�e��V� �|�:�����I?��>�i'�uXֲ�ͩ�
\0a�6����2-�*p\�a�,��РP�}ho��ޒct��I �d�>o�sz�7��
pQ�_�먤�ms��خ���+��U\���kX�����r\��	!��a�p  8�	]�5�ۤ���x�x^G2����H� O���@g25�l����8o�a���ּ��`��~?x0 ��;�q�G)�Jimt��Y���䇮���mr�)���LR���p���7M39S���L�y�i/e��"Z�%×�f�^�vn��Vg�  �,�:m�C�b.��V������_"y�D���`��5V;���5e̓�3�XW�:��ډ�������z-���8Ɤf/��1�3i��>z�C��T���  �7m�A�饳<0jڨ�=�hkc�=j�+z��Y$3�~�_=q�����H�2!|�c#�z��[��@23�ժ~&�rnҘ�f-hЈ����m/њoR�R����F p�(-�u�����~̪��V[��O%���8c;���ĭ�>wCϯ���pC�;r�n�������h������mՏ����������K�������5]�S���4�ּY�r�y��)cG�W��O4!��YV^��s 8�>ܲ2p@lb}�+*�)+!=��V�Q���O�����_�s�qSG�<@�Q��M�u����8����xaź���z���٧���BgAs�^��PX��֤�ӟ��k���Ђ�K�;��S��v7���uLG?�v���R  8����44�J�5���x����Ҵg��z���X�>X9�d�Z�~���ԝ#�+��h�1�[�k�L�|ӱ�|������c3���#j��W2��j�[���~ =�=ɴ����9K��#.��D��S���՚6�m�-�k��Eǰ  ��O"�/e���Ⴏ��*�}�~D�z>{����>��'I%��j.-A��L������B}�5���f�G��*�p�����|GNu'ň4�N']�/�4�u,�?�~1��  ���2��c���6T_�U�I�U��+�A����dN$c�V�vR���?�/d���   ���;�2�WE�	<��>�_t��:��Y�F��ϕa�gk��oK�哎E��A�*OQ�W���s@tl��S���$��s��X��;g��7��i~�I��)7d"��7��M���]��p��3N9�!��Y88 ���i��h||:��m���JQ�gG-//���Y�  y�
࿋��w�%t�5�z�M�VP�zL�����
�.�㪦�J��c����~��O�.^�Qn�  ZX�pn�2�y�m0Qm��h)�H�EJuc��
�JG՚%'.�&�}��X�r�(���a��ا��   V#_WU8b�ݓO�a��-��w��)i�^;j�   1-���   88  �!�    �@p �F��S����\܆'����ױ ��.�����ei�E�w#�f  �@p   B�  (  @��   
�   P 8  �!�    �@p<���a��pj-^�! ��!���SQ��.��]H  �8���R��h�zc � Z����n���`G�i�{O�]���   h�
����`�	 ��  �@p   B�  (  @��   
�gq�2�`�jGJ�mE	�W�  �\�L�t�%���i���?�)�7�.�qz�!��sX�  ��cY��+?�$:�~M�   
�   P 8  �!�  �?"��O1���T5!��+y=����D�j�5I�F�ǈ4  8ol~���#�O�#���ښ�V��oҽOO9�2���'�'�x6;��E8|w+��X{Aӓ��w��\��Cn��B��f~�'�3�eegi��}��Z7��ΐF   Q��i;y�嘡�h����u�ynX�]�To�#��S��67�'���V����S/�M_�!͢�|��߄�����h��ռaO\����7��:�7e���MU�9��Z����?��ّ5u����qj5r  �M�T��d/{"��E��*����`���	���֛��v�����}SQ���/-����}��/-��w�uÌ�34:m4n����m��]�7k��p_�;}�K�ҙV%�&m� �����lvT^�p��u�����ݓƬ��d�ʢ�R�=�r�V��^��򟂝9�m���5O�p�pK�j��5^��M��;�f��5N_�N=q���-�B�5i_  (����ګ�.��0��`ւ��c�Ԝ𡠒7�*|����a�_��O���9
���Z�4e�;������vت�ϟ��ƾ~�셋㞾)o��2�   i��"7oF��ƾ�˙>2O���Aq��伯-��7W���Ǻ��?���v�vw+�N/�MU���"���H��()��Lk��
  V�u{�8�=�^瘣��n�8�fL������G���\��;�|�Ls��|�7v���e��K�#�N�����g�6I~!  4�!�sÒ��#���9+;=������S��:�v���䯯\X��R��=�A� /���$��yܬ  V�q,׵J�^�m�x���^8��
�T!�Q��}�NQ��d�}�	  ���|���e�6Q$ꐬ�.��a�ܜ��93�u��G}s*q/�ī��L�k�WZ��˗�+�`�	  "}y�����Բd�K�<���lX����i�*٦l��Y~h_UG�EjK�nN�O�oZ���ZO�.~�  @��[���r\K�r\G˩T��Y��Z��V�k�.S|k�b?�a�,��  @#h�@���Z��W�먤�ms��H_���lX�R��dbUkn�ߖ���Z�mԂ�|"mݺ-���E  �1Z6��}9�/�I&V�g�+O��
��$�L����쑆%9���=����C�%sx��9χ]�c�nD&  IA{1˒��|o$�a��)�e��3��vT8��𛦎����[H&l�x�����H��Ɨ�v�^�u� ��K�h��	l���"�N�W�U/ߢbm�zk֔�sg,�]W�:��I#:���If���GM7w���a��m䤑�{�M�  @z�M3i�{f-�ܘ׏�<��^�l��5z�MϕM��׳�	U&d�|ldR_}��$^+�R�F�Z�_o���~Kf��Ր��85�}�f�I�cKQ  �۬�����~_=��ᆼv�������R4Y�
��q���es��K����p�����h���tq!����:�����7�׌�r���:]n���V�   �t��x�7q�v��q�nl2n��[�X��G'�1^é���ڵ//[S��Yo<������<�;	��z.*ۛ����_aJ�,�	?�q<j{�QG]�J�}����[���   �D^����$��	;
�·�^�}�rc&���ռ�Mg�z>6���c���;M�����v}�~K�9��Y�~�ŶR�JV������܋#�4���$ӊ>���*����D�(�>D�'BF���e'4  �PX����G:��=w����>���O�$Z�*=IжN���iV���̀��k�LiSV�v���0ߑT�S��jY��tt���H   M�U����eg�<�Q�9^��v`/m   B�  (  @��   
�   P ~���5��앫\N   
���(p(�ݓO�a��-�5p ��SڒY�����&��_o9��Q��a_��^NJN�\8G�[w�|��N����g�)�2�)a_{_�q*�W�U��>W�^oڳ��Ow|Kp� � fL��v��M�����~�v;�-�֒���;8'��?�LI��.Ki*U�"`?�;=���g�BS��R,�g�~�'* �X@DE�,�lO����y�,�l��lf������)3��$�{��}
�z�T����*���`�՚��7��^�ih�1G�w����o]�$,�a��}�q��l�a���	xz!'� ��<���p�5W�}��`kR�v�40�S/ȷe'�gͮ���*q��r$d��+�c3����'w��5~� <�H�iGJh�ɚ�w~��*8t�W0
�b6��_S2�ZX��`��K������*�_����e��n������}-\���[�<�	�?v�������.�@�2�8��pBף�3���@My��3Ϻ�vM8��G��������EYyq��8F"�wH|�I���J8婛�n��m��۾�E#��`��w�k�* 3���ɜ�w�QJ��{_x����G�7��c�=�&�YY�l�4BNA	xS檂�<ox�]%���;�"d*�-s�yZm��K��i8�,��Fܾ������5����G{��W�]�?�2 A�A��`�ɂ͟6��������'%?Ö��'���%�[T����� +$�&~��W���*�vQ �O���ǞY�����0��%"$�A����ADBNA	8AAd $�A����ADBNA	8AAd $�A����ADBN-߮t��/�>޽;n���
i'�mK�
t̸1���1�M����p�?�������O��ꭉ� �$����y�[#�D���p���;tk����uu�FۉN~$���s^��D�� L�� � 2p�ha^^�|�u]�}�|��۟�r	�۳��Մ��Z Q���Ac���5��]�\�7��BQ7��c0E��{C���Ч�H��n8��D�:�>O5%�{8�a���j�^c��ᒉ������j���}��AN-�GۿNy��?�Iy����,�1��iyJ�[s��Kף�`��]�dxܵ�*0�~�ɜ�l�v��:��`�����;�Yg�	��#p��<���ADBND��鯖�[��``��ה�]��7<���`&�����%����Mp�e|�M��[�/~�dv0�G��^H�	�h5�ڱ��*���~�����ο��vk�~� Z/�����gީ�#Z�>c��)
�S��U��]��׼� "x��HN�csB'��� "p`�Z��� N�����KU��b����҆#4��$�` d�9�E��k����W�A�� AA�J/��9�`�3��@����B��E}��!�.��e�~e)�?AD�������9�`���5I2J�à��l�C�ȁ���
OA��$JpmQ7($�T2R��t�?�I��g�m^ADc��9����`3���Z�hG��Z�;�~� � ��C������������8�r-� -�K���\�մʀ��q�����������~�l65g�6����$� ~��[��xs��w���KU���TZ��j�+�u=�Z[t���ף���[�����x
{u��i�:���GҀt.���u��R]sZ�Z9�?��'̘ ����/M�mwv�7F�n�_^�?�+P�A	J�E]!˚����޷��e����\P�RЈW؊岿v��'!9!M`��-�U�n<P��Wϯ| �Z��;�9��:�����G���?��m�T� 5k<=Z��k+�yc΢���� ��ۄ���:ԑ�PV��H{u��:W%ADL�cs��^�����շ.�w�c��Y9�e40��m��q3�f��hn��T���Ue7�z��碷Ŝ��|��g�I�׌��]�E�7K�^��jk]��,���p�����:u�!�����bLw�yy��kw%��
'�  ��X�6ģL���]���3��������E3�)cW��?�����-{�+�ʏ[;oٖX�����{�;��sFe[;|�k�M]��~�P[���s'ݺh��%_����O��]b��|�"���f��v|͉`�WQg�yr�Np6}r ��j�v��_����|v� ��`�#
y1�6��6T�ƽ�q��pΒ�,S.�|xN�kf�Ui�����x�$\X>��5S.xrdn��̼���ޚ��M=~����L��a�y��>̙ۢ>�k_�h��0z��пcO&��
|�w;,��xs�
�~�/@A��	Yyq�m�T������5u��,�O��_u�3�L0���Ǘ�]�.�>���Y|˾/���h3֒�p�a�������(��������Q�,�,�v7z��G����
c���q/���G�ی���[?�)�����Ӡ� ��Ϗ�e��V��J�U�:�sty�Pkw�dq�x��*w?~�m��ר�/�ڕӼ�>Ό������{?,Ou�O��ͻg�z]�O�ކ����W�m����U�N)�<]��2`	E��ڝ�D����]|��p��������N�� �`S[����^����-M���҇��u�{Μ`{��gA�몆
�T��;S�\����Pd�uwb�mł�6֣,�n6��ݾ�y3,��s�r�w�˽Vb-#��_�N�Eз���s �?h8�<{6�sÃ0tΕ�Á_� �HԂxT��f��P@Em3E�+5�y#��b�xy ����>�fRzڗ��X�Sd-�.�^'�_���m.�o��wW��Z������k̿t
s�;���3�N����� ��I�r �Ƭ���`��E�'F�5�r�g�wϛ}U�f�R�pX��I�R�O񶉖���;�,PA�����y�<Z�>t���98��;�}�m���ADr	�å��mf�G欦����LZ`HD	��7�+YM�=��V3��^ �����ftԑ��=�k�)�w�
wܳd>���Yu� '�H%�xss���l�y�*�4c��Xf̘ Ό�C�<�q�9&ɷ�Y��w�1��o[��A:�*��i�6�{��|�7u�;�A�<����1t
&	�$��1�E����$�����5$���0�|��H��ߌ�r9�x�*>H�z���[k��k����9}�b%��m���Pq��J����M`� �ࠬ�ݖ'0y������E`y���k���X0�n�}ȘcKg��?b��+/Ō@�Jo���D��,e��vr�A��'S���^�'s{C�HLW�k��cU���eϤ<f�N}����c���v%	8A�����-�ƪ��E���Z�r�ʔ�XN�qDVw�n�����ר�_<����DG�^)�
8�$�q���*�K1�o�ւ���d�n�P���`�;��5L!����ꞯ�8AaԂm^7��7,��^�.�v��oH�����i�O�${�œ�Mys�9��Kx�Q���k��1Lf�=w��S.|�9o
������0Й�z�ZW�����N8�Cw����mO_���iZ@�G�g/���CV��-� �h�\1�Ⱦn��1/,���I)�㧌=k�#�4�y�ά�U�ƾ�Ѭ%;��W�O����C��.�%�������}�2��w�,�I0nڸ^���J�U�
|��:��v�+��g��f���w������o�w���r����
���s�O������A�YQ�0^E��^M8ks�� �KɛE�BI'd�Y;G��FW5��W!7FNx���;s?�L�0`ɬq�2�'�0��\��1�I�wn(�rn�Ms��\G�)ΧL:g�i���u1��y,�uq���?�+���c.�2f�1��7�Eޯ*M��<��J������W�v!����m��A��@�kl�פ��q�Ĳ�����kl«hw��h}jo%�PP>еabAǘ�;	6��O֩c',��d��1/�v���sd�`��<�^�3O���Y�����Y� ��މ����:���E�L�ɭ�b�������:�3q�~�s��YK�����)��,X?ڞ�ߚ��N��kS.��$lX�J�>x�Mp�Q�7�ޘ`G�d��p����uNa�j�I�|�*ŮR(���|Ѣ�wO�n���ۢ9KcF�_pǅ�uu�)e���0��*����w�������]2�WV�EJ��\��tS���˳BzJ�����#�o�~���Tu�W���uh'����8�x^��}�tO�;�E�i�V8�ћ�:�ECF��d}��6hX�T���&�8ظ۔:7ADԆ�v�]�z��7DlH2 r>t�e�C����� �p6��}��w-���՛	4���)8sH��3wM�RY%�[4�v�=-�?`�xk�H�$��K�+��@ ^8�*2�p�ow��8��*�]�ۃC�X�9�W�k�%{X��%�XOp� ��(Q|�V�닻�6��@ñ�	zԜ���gN667?o�5��\�x�l|海���e�7� �e��S/�Wua���d��Wj*�P�~��^U� ��m��]�%*\]�5fdz���W�A�_�*aa���(b� �H��^�޻�t������xF	8��7{����R�-��Tj[��&��{���N������;��И;+K� "���k�J�^�����W��9�Vo���?�rEa�l�곥��5�5�i��e5A�A�������Ya�#�ڜ�I�A;^Ǳa����Vk��O)�7� ��ڥ/���i�qe�n�v���v�u,�������o�3_?�hh ~U[�n���*=#��ߪ-p� ���V�=��?��Y2p��hvH�	� "!'� ��� � 2p� ��@H�	� "!o�8%;���GܟD�*A��!7lz�s`�qg@��G@��Շ`�֍���%I54y���0��3��N�����2 "��U����z|nlN�Ǻ5���j�{ Bn�9�������>;u�y����p���u���5�=�r���窄�߭����G����g��� ~�l>���k���)D"H�M�.H��͏ÀN��Ƣu~ŉ�ax�c���S`����^��Z�sN!{\��N���6���ؼ$�� �i����=���'�?����C(�.�.����!#�Ǟl[����ɭO��'n�/~�A�H�S$K���]X���Uᯯ?��p��=K��e�΅G&��Yy�kςnz�=}'|��: � �d!O�}�e��l�������w�W�.�U�7���c��eQ�Kn���
K��� "H�Sdh���?��MP�;�Y~ N}�zXx��p����&���us����>� �0
	x�`�y��w����.���vX���0f� ������g�_/� �0	x�`z��3t�W���S�?W�.2
+�?�D��\��oA��j������=<�C  M����������j����XK^��������M�U ��!O�JOM���<�zp�����%�M�����x�9�����f)�(��o(�$z�}��j�����l6���}�q?n��SEQ!��~���⚊��l�`�? �5�ߜ���K��Ώ�
�O� ��	�E O��%�{p�>I���z��/���\�+O�rş��T�Vo	vT����ioY��E �V6
%�Y�
6
�_G+�1AUu��t��B�a4����$��n����	�'
|hr���Bg�]�9�"D�����ȲA��Y�����G�'W�����~�+�@�T��0�wB��
������uѶ0A�Z��Oanj��]�^�.��So�$�ZG��t���`��ܳ��L\}�񍹷Qtm�p��'N��4U�-z�����1ץ��2^��ic㫚���~[�(��ص����Ǳ�h>H�Sd��`wE	t�/��N�|G6T�k p�����ek�7���~�����|P�����(�.����qmE's~=�a+V�x���`х�a7��m6�}g��Eԣ�g�ZT]h}^���^w0�-�E�Q�u���� �[s����	[��	����}�u�
��DsA�"�C�����o#'����N��&�s�A�i����D���~�G+�dK �0�U��u������-q��QDm�.^o}�phyot�E�Ǿsa�f�0���EL,г/뢯����".�wp�h6H�M୍�0G�8�2x�������,L��xj}n�z�@d>������v T�\�2Z�\�G77�K�!w8��rx��]��܌�3�{��\� 7���ќ��� VX:�ʺ�\�۱���iش{s�#��{�8��]@q3[��2G׸q�\���Y����7Z��u��G@x2���A4$�&�k�F��$ÂTԥ-��b�5�`��0�C/L*y�(����(�h��!�8��OKȓ�2��0j�E����F �	��D3�R�C����x�	�yk0b'�M��}^Nk0���-a�&o����&#,
^��Y��'��v?%�D�BN�{�ӭP�p��1-+*������YV�%	-�t+' �6�p�k
(r��fQ�Y����%�������^�	'�愿����jq杪:r����5��_�2U��>/l�a��T���D�20�(�H4&�h}�����#��֭�fԂ�\q����c`�Y2�7
�Ȫ�Y��A�5.�x*�n����[��*�Y������	}�[g��xDL����p �Dy�8^����Xx�Ğ8BXA��l8G��g��\�����U����@��-k�b��`no,�*I�Y<{�����8���Qw6
/��c�7�nw��oc��.��ذ:Ad�xN�)�aY�u��
။~!�p���Ȝv0<� V�"�^U)Ȕ�B�bc���9�0��o\=/˯��f{�J�JgQ�m��%^�(�l\W�'�:w<��L��jp��O5�V�d�༼�0J���X�I�Q?�r�`�#�;��)��\D�@18���X��$���FcibXQ�cNw��@8m,�O~}��G� 
7^SS�����XF�v�E~MQW($�T2R���?�SOx�d'l��� Z+�z�
����aIU�Ür���D<2b�T�jRj�k������:�EWܵ>��T"����M�f��e�u��� ��hGln,���쀟�n �ֈO�prXg���֛ڽ-\c��v�2�2�נ�k��jl�x����Q�1���~�0ЍUz�3��+A�&���]��o����U�c���۠�pzq�U��+wk�*�:ج��"^,Ȳ
	?iA�A��}w��wTj�#Z��F��������7p��}b���5q_�p�QB]��R\��M����I��|� 7w7$޵���C>��* ����	R���[T����r�"������)/��^�e��.�����K�ҹ����up���������1�/��_��&��ǖ�)�Y�./�[�e�������;ם��9�F��o��Ǭ��u�x������&l6����F-D�V
~W��5 ��c�ϵw�⻷�/~�̕�f�fL>���6�Ԟ6g�	L���]�͆����}n��J9�B�@`�������λ挼vO�ͅf¥i����io�^4'�>��i�M�{�ߏ��<�m�=�u���\XWK����e�y�n-�H[���nj�4<�)�mMKMlEQ`���Jo����M�RNp�Co�3��jM�][u˛s?o����O�M�2n�Ь�8��f�vKU��qu�u�?����m1zռ���M:w��_w�渨JMQ���=��9�>1ẑ{>�|�W�9ۭ*�:�1�W_����ch�(�������u<:�B�#����zT��aw�A�����q�Vx��/`���h��<
t�G��f�UJ��1x�k�z
p*�Up���3��Qm�u������̇TY^[[q�ҹK��9���N�������|�$��򹽟U�Y��Ҙ�6�Z�k�-ے;鼑9���F֠�s��vW]�Μņ�;�;s���rǅ��[�ڹ�3�"^����F�t�?d:��w���b�p�6ֳ�3��3���?�kv|�x�y�`˗@�M��]�X�M]̱�Z�͟�K��v{��`�X��Nf<�u��%Sq�A�M�f9������Ѵ�FO�Ɉw�w���0yܟN����h1wi�=���k~?n���.���U���8=��&3/�[w��o�Z��������˝~�'d�O���xgn����΂����1����a�M����>��_�	�>m�qyA����c7v��p��� �T`�d�`R�^ �2��1h�ěh�s�������g-Y�Աߚ��9�/�jhV�Y`"j��x������7w�;�����k;�6���{�՗�:N�U��B�����鏲g1����Gϱ9�;���;����ϥ{�Kݢ�vp7�,�.�dMa�����l��t���ݘpw���HX~K{8m��ࣲ�m,m�)]h�:8���������(��An�t��� �)���,j��[G@T.8z�,�����U
Z#Z9��rUV*x�5������c�]-���,{d���9�nkl�F|�DЮ��]��x3.l���݇�~X��8Kg.uw����������Y��(�^9=��pK�xc!���/��?y~8�kR���n9�����؏������;��m��R�H����	��,�`KР�ݸh�b*�`?�Ǝ����7�.��0�M���w�X�x�@g]�l���[z�Ҕ�,}xiY׻'l�� &�_����2/W���w�x��{L�үa�����bZ�cn�.���c�~���u+�ܶ�Ic}�g\��{��M��[��eV�_G\���ɕ�vaJM���z.>N&8-v�����n�H�8� �"�)d��H�qVm�Bø��O�ֈL�}�R���Y�)��o�w��!�����	x[�'��fx�|`Y&�hr�H�kz�̍|XC?���y���ɒ͟����w�Z�]��a���@�MPPq-;��b�7�L�BL�!(��Ȋ��o�[�F1�m����qK�����	��_kKT`Ǫ��Y�l!2�DZ�rӢ�� �t\,��_�"~��}�������f_�ŪϘ,~�L�+�m��M���%F��ymm�� �c��#��:�6����+h��jܖ�Y�v&�, k�'��ƴ/�nsJuk�^������8�����$�'^7F��5N�^���be�v�Σ,�h�O��?2i�!��!��s%����~�j�@�V�K�)��M���h�3����w��dJ��	`�;����5>����Q\���l�ݦWr��,��1�ǓtQV]��p|��^�P���x�!�[��h�(	�����S��l�y�*�4cI��3&�3�����갟r�I�-pLz�Д�4o[��� ��Т�G���K�^S��U���9jR��#Z辎o#Qݘvv}cĸ��^O'(�\#y��ҫXqK���Κ�x��	�:���_���S\ǘ1�Ϳq{N�6�F7$�9"�r�}���X��ߌ��ҥ񶕨�@��4�i��u�?M����Sܷ��D�EO�Z6*��<�Y�d�<��1PMN�ۍ�c�u�ƮK����M(��Q�ğ\�	"�4�`�y
��E`y���k��w��c�$���c����4�T������X�|?����[��J}��f7��=�*/��x�ɥ1ђ�������c�Kk+a���������1�ިxc�5G�hZta�&Q�v����k�
�`���㫫�,���p���O�}�%�X�ҺH���aVtӒd�p㈬n�c0�D�`?��~�
�œϟ��f�"l�>]o��(��SGT�'�91�Pm��X��tP�uÜe/�|mt)>|��p�г���o�{߭�2]���!��t*K�|�03���Z��Њ�̩4b�"(Ԓ��W]�(����������D��P�5�X�s�y�J��D��`��;��ް�K{A�:��a����r{���ͬ��M��^4m�Էf-��h��~���tN�`˞p���/���I�Q㧎=q�3��x�׹���Y���e8�G?8�p���q{�Uض���UeP����9+��W���ԋf��W��ӫ�v�h�H�՚`��cR�r�h-��7��ƥ�7�)��I4������J''Z#�tC*��#�����|ދ�g�)c��<��A�,S�Կ.���ɣ__>��_��W�O���Ń����fh)��!��w�Iㇾ;o�w�;���}��rVd�i�R�)i���Ѽ>s�w#��&D��iߕݒK��^����)u�"Z� a�8��Л�"�������.dۃAmhcw���l<���D��iccsv	<o��xh؂Q��� :��;K�.6��`���b�c��A��ܴq��Z�T*��)cqf-�7CK�B^�۲7�'��wͼ�b�����0|�Y���[�ns�E�I:���(M���g-6Tg���/>V��O� ���YVQ�6�y$(�X�t��Ep�9���cF@;gnRc`D��W��
�� Ѷ@73��]w<��MM�5��ʘ�-�?���b���-X��Y�*����ꮑ�w��"��-���8�����;�i$�D�5���R�خc��E�!r��)c&�=g�"#c^4y��:s�o�V�H/�3W⬿Z�8{��?lн�����w��n��ނt��3�5Z,�?*����x�>U�u�����o���gu��<ڑՏ���_}���Zt�������̅�z��<��d�O�ǲ��j�vW��Hv,����-��nz�׉�-�~���%i]���Iխkv��"�-��1�ъEV�~C�\�~U�ԪOƔ���7)/򇻥���pJ�n;�G��0(��H'Z!�j���yHs{;^F�_X|��-�-�,�(�~�u��N�����0��n@�f�(��#�\�⫃�S�<�jmx��+�g�X�:ЯP�r9�q����D��#�O?�����'�L��x�-����B4hl�.|/��n5Q��#���o؍ ��R�j�cC���<ؑL�i��.
1�ΕP7g�j�����mce7�~Ѕ'�3�>a��!�A�I�����)�<�%����c���M�@���7 �?��|�4u�ϯ����\Q�(vх>��M �whn��Cr��9�SU���A	v�8�D�G+�wW(��~�j6IU������R��I����P����mu�e�qk�Ͷ9$�j�/�FĻ��h���`�������tڂMXX�Z�NN�bJ<{p'�P��F���EIjR/�a/h%��6������&^'���G3��Bॲݰ�Sњ��Nm�p/�hpm9� F�>y=�+��`�t�'�c�B3�B��wR��(�r���}k��s��3za��{�9���Rs��ؽW7�N�?	2��.x�t7\UԵQo�d��W�
<��!~��Ε �=��xPj6
fS2!����WX���-1�K����]�(����O��\�E�<�X�'yU���m���@��&w5<V��.�32=S��+�߅/]��� ��1C�^�ʶ�Vv�k׮1-����SR)���n�o$z�x)k�Ǎ(�	�{��	��c����]�`�A�B~�"\�����p�>�Dc<�S0����R�+���9A4\�F�5R����2�Os���HP�R�)��Y4��f�@���?l��v�!W���&'"��Ƿl�-qw��,q��R���J������[�9�Vo���ۯB���^�[�.��]��F7�Hv�^T8J�x�z|�Պ�rd�b��1�͎p��1�;����~�������u}.�]��:��&�D�f��Jw��j���l�ksBg�� v�ʂ�Z#�Q��*�՟�R�o$�d0R;:%��QENP!B�U��m�Ni���-�<��0��}�Ǹ5�9P�2"p�Ե�����p++��3��y ���'�LF��_�G���#�ڸݬҹR�8�,��u�Xu��H���$�a>$�a2�:Z��c�,2V-�7�L��h5Q�#�3ބ;�1W:V��l]� � '�������l\����l\��k���#�2Q)I|ߢ��H�	�tH�	�d���cj�g�(\{nX	ע}Z�9��Q��׬�>��Բ���@�YH�	�d��'ʅ�@�$7��� XA��j�G��Ds-��	A�Bn2�g=t���>�m�ĺ�%�mg�N<b {|�ks��]D�'�E�@0#�G�7>ME`Yq���M��I�B�Edڛ%A���5}<?��o��(s��	v	rrsR3<�WɼJlmp��i��n�|Gv�m�*���|���P�'{{|����'����G[�<�\�M���na���h��K_mbU6������<l��k@��?|^�E�0 �1Oz�o@�,$�&��=��+�n֣|z���G����O�Ji�$�J�{d7|=�'�(
MpA���#��p��/��|<lR���`��8^��P� )8A�
	�	�pJ��Y~ J�ˡK~{�[�^�������?}��l�$�9�q1s�c��kX����%uNo��x�b;��#��fU����s��Uh����WS�&:A�	�	�wC��e����[�U~Rρ�B��X���O�e7��<1	��. ��.fB�:1���R�8���X�"�t&0�{��hU�ހ@p���C��à c`�/N����ĵ�x�hX�5��G4=Q5*�BfC�"�v;u��Wyj�G��D<�5�|���p��	0�⛁�-�὏��oy�}�(wU�v���H�y^ц�<��Ux�5����ȣ�E��-��7Z�(��
�`�rCW{�8t�~cu�u�BMOpHv}�HT6	�r&�>��ʴdDfC�"��T����o6�0����'o���w�[�́\{߽,��_p�����X{�h�i,L�w��E���wc�������q�5��jC���{|�
��~����� ;�YCQ�x-��~����d$rM=L|��HF�C�"=;�=^�������up�.��B/p��1]�[��3����m,��"�ӰQIXd�>x2pqҵP��X ɾ۸?��t8l�{:>��a�F����#���� ̇<EВ�9�FX�ss�t��P��:��Oo}
��_�WUD惮ot-GZ��-{e��=nRe2�;y�w�n�;�l���%B�-wE>�f��Xpg��~}��{��Y� �Ð��Hd�l���qX��y���7�:��Q��w<˄=���,�8��j"x'�G��u��*��6v>	7���	�ό�,d]d�������D�c��O��>Y���c6���D�A�"{+�=>�]'ذ�'���x`'�z�F��5�z���uAG'2�hWz�����N�-YlE*��S)�	��_��xV��O0">^5�ÉDdN;k)J�s�hVH�S�=��cd�[?I��mw�ȇod���:���`�mO�Zo`d�]��Y��X�<�������Z���bu׉�?ņ׉��^���򮸶o���MQ等	�FB�v�x��w���6�1��؟�c������C�"+�m`nt� �ECF���Mؼ"������V���*��t!�����Ӳ�+��Ha��v�0�L�����[%�+��c��L���ݺ����Cv{���f���J:'b�_o~���	x�@�"5^7|��Z3�TVu�#���*�qv�`�t��{u��B]��HS)�"�5q���D�O��K�R�5�h~H�M ��(���s/o��#�+J`�C׳/�;��m���j�`j��˂�"�x�������a`Zr~,<A43$�&���U0��Euϋs
��Ӎ�hg��&x�wB��j��Ԯ/���`L��p���"g�J�c�n9�/�;���ڑy�>�O2�+�j���"��� �BŞ�f�"��N����E�YuNf���z�D���#	�uE�_�&�~�P��B�s�H$����	D�Zs��^I��yՑ�e8!0#U�̈́#ȱ�iS�~��732� �Đ�D��Lx|����|kL�
����,k�]��lC���M���I#'��ANi ה�j�5$t��ִ���pt�cC�To*X5l=���)�G4f��� �	8A�	�����$$/�~,s_L3��-�`?��>�ML��lR�x��!"=�r�K6Z�y���\hid�Ѭ�XRأxa���z]�P~
�����"_g��=�Y�l3��Eܙ%��p#�U1`��E�����G�;g��������eA�:�vh� �)�����_�S��C8^���Xx��X���bA�~�,8;�ܺ�������eL�	"��t0���P���~�K�۔b�:Vz���`��vl���5ir�DB��NT*�Bd(���iÜy`������E��A8�v��!��] �T�w���"s�`6�.�]�Е�iX������~��u�q'm�䖣x�{�cYW��j�f�lY����ǅ=:��NRe���ؽ��ܸ����b�[�kc+�\�$�<�U��:3�:���]�ON�jA� ��b���G1� 7�ח��
/6�?Y��Ac��P��ҏ�w�Ne@�b��V��6C&�Y���Eݠ���d���H���I{���]�7��:�.p�E/l�"<����l�]����FÛ�-kѐ����x`�&���-t.��m�8&θ�]k{}�ޤ-o7��I����(��+��,�L&�����?ĿJ~��^D��.sL۲�=�5�B͇�Ã�h�u���~Mc�ߍ�����>��y"��5m��1B"�k���uLg�zeӛ�Dss����w1���w��B��)�b�g���/��W�%�|���Wa������]6F�$ #�\����*)��� 0��U�e���ut���`mNV���sA�Y����T,�$#ᣛ�D�����xq�A������o�q���"����軒8.�X�99�E������;����h�K#٫�L�s�%�4��4�Oc��v����{���f.�3b��Pν��d�����%�eeYy���<V���㈌���Eo�&
�c������12�Y�q��Eߣ��h"A��38}�u���ݳW��,*_Z9se��	3&�Y�������(�4����U�i������_�&@pm��/������w���\yF^ѳE�Ԭ.v��׻*��1k���	}���m´�=֑�X�U�9�ks��<X���D0B]S4��ֱ,�n��hҋk�^�B�r"�9���u��Z�_�T�����O��'d`>���S�M�̛�O���=���U�������-�@�z胗���|yZ^��n���@�����U~�9KW=f���Ox&�Y;,+��v���^~{X�?�����<8���WQg�q>�	��V�}�wxS[��M�h�Q���ǂ���O�3t�3�������}�}ɯ@4���5VlE�c�cP�1�y[�Z%�:��M��N�L;/�}��e�,ot���h�_�ً��SƬ>>���<��,��n����Pِ��~�S��qO���?:&�{Z�U�27���T|-������0K�.]'L{�)�v��c�|�x���}㮆�fT��`Ƙk��^��n,��՚_����<�}v<<����� �_���c;v�G:�=~��e$�)��.��eY���X�]�Ǘ����2��x��v^}�ߤ�d���kB�8�bnMltՌMF�à�M���΂׍��'C�*��֔�O������s��+�6���7�yaߺk�_8��M=~�%�r�p�0g��Xۏ�-ޖ�g�|�=0f��Udxs�
X���i�6��`�7�`@�0v�p7�4���²ￄ?��PVKK Dg\�F+Y��z�D12ܡ�/
��w:F��lB]:�+
�c��]N�)N�5!�]կ/���æ������˽�⫇:s��5�+�`C�}5���o�+��΢�n�E�:�^��O��s���*W���ؠ����ˤ%��Gw�%7>}�w��L��]Q�`?t��������cn!��g����a�]/��'og�"�in����ƨu|�nn����L���%I��6�I@��\���g˂J�e�,XC��cQ���]B�թ�c/W��#5gicS�Ǔ=�����~�
�̙�b�w�.��͸�����g~���ҙK��OX_�%��k�v%�Chz�Ŧ�B��͏CQv>\��,xa�C��*��^���^��nX~˿`��Wî�@���x�n��z��0��X��s�嶲������(t���Z��9��K�ò��`���\:	�⸷w��kW��f�B����	�t�ث��h�5��^����L�
E~L�*���ߝk[!�.�,���W=3}���>���r��u~�sÃp�w�'!D�S��xd=�0�Vn�'� �R/Q�=]N�Z��xw�'���;�7�����q���q����Y����;S�\�?od?Cޫ=�" ��!HXփI(��e�m���v����	p|�~pϒ�M�0���.~
��W��?�}��G׹$��M�����'StyK)ވ��`���;����K�D��@�q5$Y� �Όqp�}�T����!d�ϼ�Wlɴ+��~��Jy��m-��\{L=�J��t/�� ��7�k_&�?��϶mLx���Gñ]��o�n��v|�>~�8�<������U)����Ա��E��1�������U���ƚ�X[=Xj�����%��|��+@���D�<������f�G	XL�6_��9s�!׫!��s%����~�j�@�V� �{D��-8n�y~�[����f��.|��{=�&��̥�a��Mpڼ��"3�}�w�,���������HD0�Kѿ�@�r�w�\w��I(	�����S�3���U��f�#�Z��{���m�iH�WdI��m�|�+���4o[m���կ��͟��(�g=��g/�Ը;���73��䞃X��P���,m��S�&��Z����1�O"
칆��U^��ݸϴI-A�)��wqs�MЯ\�[PCLpQc�8�8�$�?Qبx�|�p�D>�O���7c�<^�,޶5}�_��86��
�`�y���m�����4ޫ��ou��JmGu���%��y`���c��tQᩁG� k� �� SZ���;�����I"�dJ��n�\QĔ��8O'\&�ˋׂY�AǀIt��'�8"k��+SJzĢ��xۉ���~�'7.�f�����a��b9��$���� ��ۮ��pj���sVf����.��^���0	�~X�P��䑈��>�˖Tc��&�NY�MK�5��d&с��7�_�>a���U�g�I`�X{A;��L����S�B�z�?y\����Z�"/@����5��X-I���Be���"��Z��/�rUA���Mo?
w�8��1(���"~�x�`'�m^�!cE�$u�<�?�>�s8�����@�&9r.�2n��sݗh�������tfO�hϾx��qg7�|��.8y�-��x�ק����M^�ux���&x��z瘮}���s沀�JO�v�A����=��`�|�ě��ڪ��r�\�:�Ņ��4)�l����td���ǜq��s���C��F����g��Џ��kǋ�wYqXyː��%ڔ��/��$� ��w��3ؖ�qV�+媜�:��A��uϷ��
��.�#������a���nG��&�w�P�zw}̃5�L�	�h[��?d�E��Q�����"L>���{I�M�*��:@����eq<7���B�c��w|7njr,.���c���,�7CK�BA�������ӏ��%���)Χ�>�����%]D{��e�K�I����q׼5w��F�?��	�f���y�eU��e�N��e3\z�9�)��U���*�d�����g�KW�#�v�Y��^�����}ŏ���0-�8���o>� �&[�߅�,����0x�88N� ��^ܿ�@5ც����N1�wm�s����ǅ���1/������Ν�������6G�P��Wq�Y�W��hE��z>v�'v�=�{	�(�bnk�X��W�R�{&޽W�LZ4{��X��������ю��8�?�����5�/z�d�*�lع0�3�+�3�Y�^�qǌ��:��i��#���~�Kès|�w�O����#���gV����\ݘł�p"@DۅY��E��n��q�cN�l�:��a�ڥ,s�0��5���M�ݗ�@��Ӆ�gL�a�O�%��Sƌ�$f=t����������,�3��O7�/���U����[�\�@W�N����c���	~ �ٽ�A��c���R��{|��ɯO"�
Bg������Ų�-ҿE#Ƨ�{<������ޟ���> �/���l�����-(�w-�|�����9�8XSoo����3V7\U�1�6���o��x���K�q*oa�[[f�7�[�`��v֌$���(�[xb��`|�T�e�T��9�����n���-��us��L�����o9V�ÿ��#�,���߳����9?[+V��r�o��Q3�3ꖊx@��X�x�xЅ��g�x'���^,�wu���	~k��s��o����2�!U٧��qX��D�s�����r�G���b��ղ����w�-�r�R?�v����d�È���?L��2e�0�m��g�˦���~u6{��a��G'��ڋ�]��|��xX��z�����b��8�M`}��:,�֙�=v��f^�����P'.V�Tk�{<��v,�?|��1CQ%�.9��v�������A�a��h��D&�
VY��l��d�}�m����jE�ĉ�'���mH��)NPd�=��:�6V�U�#�� [�Fm�1�X�۩��w��E6���N�u^����8�ɔ��h�?�����{ge	�sP����]pc���7�%���-i=jNp�|DvN��p�LPK7��������C�F_Z�.r:���Á�����)lN���K`x�c`x�cX�8��`pV`� 7\3s㈋Xc�?��gV-"yPP����5
�M���6@���_V�Ӆ����NB� [T��!���	8�*G���
54��X��eg
%��'N&��'�(���[���
Nj��G�[�J�#Z��-K�._����Ɉ �q���N�q2�r՟|������'	�	F�oz�)�v�A����e��+��`i~xs��^�)���ݰ���V*�'>7V��,̻�f�^�n]�OY�EX>��5����γ.���n�e����M��-&�"�?���XLZ�(�h�iP_��(�����5����N��Ï��<�3R Q�%���+��9���Fq���u~?�
����k��N^��hy�-z�g��OT���=�_������?>��fb��Sw�5E]!�O�G�42R�q=sMm%,ҿ�V�Y	��g>z,��~����,=쎷g�ql�#��o�ӏ
�vn�qO�I�L���:5��~c�-
R2��#��M���ޠŉ�h�2����p�����N\�k��?+�-3Կn-$�Lt�����S0�Q����ۂX�E��7�W/�Ǔx7����}�a|A8љ�4�3J��]���
>�*��r�j�'CIu9�z�Fx袿�_N��������T߸{+�*e?�X2up�>�Y	�K�װi�mo>j�~:U��bZ�[�az�J��u!��(.�n%��7��,u���m���v����Ѱ(\�Z���!j��oIo����b-K`�_����s.Ư$s��&���pMk���b۟t���]��0�_�W���'Շ���B���(�z�pL��V��S���[߹kY�ykǧ*p�����>}��{�4N�90�U�Zx}�G0���`��@�0X���Y�����R�}r�OЅ��^]���h�R/�]ӿ��� �x�e��(L��g�(����8�����~dPp�v��Ykj��x�/'M�^��4��߶C��p��hB֖ث���A��vn?pdA_[tlXLl���o��ο�j��]��/e�F�2?��+^���>��г�3�����%5�l��K�:�'�A	\!h�cdr�ԣ�OR��Z.Z�^��^�Y�&&F��
ԭ����(�Z�ڃ��<�aڕW;lͣP�Z������>�}���|�E#�#	?��3�l2�od�c0z'�)��Df���*vku���P�Q�< �Vk��%0#��F���10-F�tS�\ho��m5�dE&&�C��*J���v��P�p��b,k(���uq2��
L���[��.�ia�����g$�'��x�aH��6Z��k�7�bc�K,�����P��� �Z������u/�B�����l�^I��q,-Kd��7�?��`n;ϖ/p�׍���`a\��1v���+O� ~ː�m���	]A�m�H�Lh��-��jc��(n
��jM�3C׀1:=\إ�u��xf���-[,�^���21�	�{1�����S���Wa�.���������WE��Z^����.�����gu��pi"����k@�	8Ѧpű��j��V�Z��f<��E�ǈe�$��X��'���yꁸ.q��v���R��\���Bٚ�o�;���ª�q�:��1���<�h����\��F�>i_��$˝h���m�D֜?F!��"!	�6q�9�el<,��WZ6�"溽�c����ʣ6R�E?��Q��I�
	8A-B*�A��ADFBNA	8AAd $�A����ADBNA	8AAd $�D���8���_i,���5TYkP��qV��Œ�X��5V�[�	���ק����`�,}�uZ�K}"XF��`ŰX�g���J�ZY/Y�b��`mt+W�<^�7���z�<;'�%g�8�װ�+~�Xߣ*+1��E�mH!�O��pMx�.�H_R���3,�*�B�}��+�m	p�̀:�u��޸?�g-(%]�P�ܵ�K������,Ut�Ǻ����c�M:P�P�,�;<jr��7$T�.���ZC�ζ)�&�������(�$�(�'���j͚R5�l�lK���[B�#�mN��ޓ����߫��4���+P���9Ԉ*s�����@�3�b������7��P����*�� '�hei!˖�9pf�tѵ6�_�������FX�2�"<F���������y]�#EP���U��き@Ђ�sE7��E�yHSAaD��I�*�|��l"��\�.���ЄH/�@�Dc���ȉz",V���G��������e�G���X�Mmp�M���Qh�}�#��EnU�M��T�M�pE��Q�	x�o��6T�"j��w���C�� w�wG^#�����k-Ч� ~���m��P8c�]����5k����~(@�Of"M�R�x|L��-St�;�g�I4sE.��3�~�g��9�����Vm�ъ%j}�A��?4�a��~D� '��h�f�%(�(lr,�.�S̽��E5��n����'����ؓDpT�.ǵ[��F��lnW1�$`�O��`�(�á_��� �..��������{�K�5�����fA�	8��rV�Ƣ�U��}�rK(иN�0�u�p��O;,��b���	0��uA�{��}�`���[��'x}�n����5���g�Y�lj��5��s
#��BN�90L3�BkS��ͬf}��o\�F��ź����xb����`9��f�r3�������:�������O-1�mv����n� �	8�%,�v�JC1S�������(��Ŝa���|���ׯ%�����Ók(�.z"�"�}r�=���^G'�y!'~�s��̊��pcQ��Þ�Vyt�V8�[�S�%*���G���r�R窶�
���F㡕͢ĵ�e��-��#��`���[��&�~�/�������o�~��>'���5�8�YDz!'~�x�2�G�[�Y��G��\G���'n��޾6{�\t�lx�}b-!��&1T'�K�v��NJ�^_�}��2K�G���B����Hp�͠��R[�I*�-L��FK�K3�~�b�\>���d�J��:YS�� 4����g�>����8�?I.;lAŽE�ֽ[���U��V������:�Vk���Z��8�u`m��m�ފ�����s-��$�@�Ϸ�!w�����g�r%�۫Mf������zo����ϣ�e5�(yy}�φ%|n�X)�iǳ�? v8ğ�Vx�!�n񤚣 '�Jy'A1�c��Uz����Y֟�� ��1�R�lc���P�:s{NZc�:}R�1��E'�(ݻ�nP�t����PM�k�VW�9pI���O�(	!��O,@S�4�)�_"/��B!{��:�}݊�v	)�����8D͓����X
��7���7�p<;~�J���B�8o���zÓJ7�K�e��0 ,~��7���'tw����#�!hh�)!��r����!�Ћ�!8DɵL�*������*T�*��Ӫ�B�U�&� F��)<V�O�� V>��9@!����\���:@�vE8u�#�yշ|��&\�'�bE}�&��-q��F�0�~
����@ ���e��t�$�ɐ��T�B���X��V�ڍ�s����]�4��3^U%���^���, �b_��^�Qצ��0�):mr�ѐ��#��u_��[%d�4�sr5�Z���p�Y��w�	��^���H�m�J��j^��;zMd��:>2�� <�	WK.���D`�e)�"�S�=��S:�E��!m{C���Y���[���kga��s:�4�4!���c�wP�,�1;��e߾��|�J���Ȣ+�����xk<^��"ɔ5�����wv�3���]sps����B�)������۴�/>�浺�Xj�*��ޘ����/Q�K,ɽ�qkٛkG������W�|���L��p,;I�&�a�9P�������|�~p#9&���WN!�����lFX�%��i�m��[��o6s��op�5l�7��v.�?Щ�2R&^�{C�}f��Ż�k���i/����/*M��'d���Y�����ټ0�C���m��z�%f�v�	�l�;F1||���z�,������?��K6����#;�qbą���7��TF�o2}l����@��'�5����qQq6�����.��:���}�;#�Ka��&7o��GO�r�es�->i²_/����*b���ļ�骍FSBNڨ��w���;N@X��n.n�"��'=�T����L�j����cf��Z��M��Îs�Yl����ۃ}��k5�A����vO�\,���}쥇��荿�q���bk�\3BS���ň���1L's��%���-�;$��|��/R��גG�^k<���j)��ի�lXz����׻|��syY;b��m)��c��q�5���.�ϙ��Q���x����7�ϟ���ص���{%�����ܿ?%셈�+aÄH���͗�x�/��Bʧ������r37�F��+ﹷ΋��1{���*����ӹ��]��cJ-�o�����ѓjK�4�A�^oH�ԍ��y���T�v�'#)qY�L��&{��j���u�s�V������eoA��`�7{<l-��ϕ��Ԇ�Iw�BHو���Uf��赺ی�+}����1��$W�j��j�r6-�{���l��7%��v����[����b+��l{��ܚ�C<U�.���B�H�t��>M�ܞ��M����-l����\��Rv�b��	[n�����T���'���*ā��D�fذĠM��:�j�/���n����+���}5�U��n��\:Q��ￔPp���B);_��>5iz��I�V��K�g5+m9Φ o�#9`��;���4 H ��A��>Qծ(����Gc0���̏����d�:�埋BH�X���t����	��6��'Scñ6�ҩ�yKL0�G��O�R�+��IU����E	�P���%݃����_�{=)˱ƵB������$=�*_ϣ3	x�6��h��|�M�>�<"��L�Gx���]HY̗N�U��(�*�7����m���1w.B!��Y���k��Y>�G��|��v�[����6�9�[��y�o��w�^�eu��/�P�S� y:7�{�3c�ЕS���1�۷Y���h�6vh;p��m�B�,0�-�c�3�� �2�v|�����J�o��Ҏ�)�]���wF<���ǹ܄�,�{���5�s4y���_`F���/V;�����>��37��?7ox��Q��H��t��?��;!���{��Z��*cIi���Hx��͝K z�
p?�t0�T�&��^���+r�ЈPI #�ln��d��rt���]k��N�D�&ܤ,�a>��h8}�2��wRs2��-O�+��o��m��N޾Q��B!����I��
du����%ёіS�"F���ZO|�ҡ�Wj���Y["w���Č��SiDE�#1�񖛟�R^`I�,u.X�.l����Ya@�h�m��zF��l�$O!�|p%���he&Ƽ�D���{��<Gc�wn�'o=��
������>�v�� ܤ�B5x�Z���D-��g��F�2����9i�(f�B�%���  �7IDAT�ᵞ#���Fq��Ys��m��|��n!���9��a6�Qk�˄ܙCWm]��\CʆM�Z�:x�t���Ӯ�1e�����~-��OF��*+r�H�V��4mX��ű����o�P�[�^g�[$�Q`q0�����B�4^�ˏ[��&ד�����|�un�7!�~��̀t�/��*�O%�n�Ma�O�X	Ks�f�m/Sn�E�/���foK��xrD���#��;�l8��ҿ�WL-��n3��r��<��A�6/�[c�cF�?�V����EŮ�$���a0��{��!�T̄�I𜗿���b���Jp^4z�¸h[�9"<��r���D��&�/U�Jt�nȦ����%j��a��q��t����^R��������j�Fͺ�˝ni���3��cğ6��4�6��&�ʦIO!��Gv*tqq����r��XO�����������~�e����Y[$���\Y_ ��K��t��߯Mf�8t���Yg�?Z�73e��M�  h�- W��.�[�o@3��A3Pmn?w�.ɠK��)�.��>��c��ZayF�K�&p��7!���cd�3b�#n�+s���R�Ҭ�v��;V���$j���~�R��ˇ���[��$B!�su��D���̪����]�����Ba�z���S,�[]�fݲ<{��f1��
� �R�=�ia����o]`JY��y٭�;{�C������+{�I�*��mj��>����!��sI�����K>u@,��=9u�'�WS�<��u4S!�ۜ�̈́en�!^۾�Y9e�c;��i��r�U;�9!�烝���A�GM�����!�oN�:�	N�d�$H�R7!��
��)��@f
�s���
7��Vw� ǰV�on�^wuyp%/����z�B!|�f����/���B��&2%Ԓ�p2�ǺDh�a����)��ZZn���ɉ��By�`�DN�9�\]<���*��F�-�W�����w-�6ξ�d�$3>*whS�1w��;p;�B!�Q�������t���΁�3�m~�֠��I�]�������!�R��x)ݠO����GwCzƩg�eÏ���k=C``�.�&Wq�B!�(��W�7]߶s����qgq�Eнa�q� �B�Q��I��o��[���Sw���]��u)�	!�An'��}���xJ9z4&e�sˏb)�[��BHa�v"��D,N>���:��B,T��7C�\u�j�����c��܅�����{���nXs��m���!��Q��IJ���n�}j������F>u
n'�����c��V����S8p����u�[v�z��~�Nܻ���Gn'߿^p{��!j�wez|H���/=,[�B��(��$��)��u e�0��hn(ٝ��6=6��&L��<w�q��	 ��^)I7�#+�%F��+�Rj�!�aP��I�&����
�t�=o!�΀nZ}\K��yr7��sdk�͑X��M��G��UJ�J3�ٻ��!!�1P��Ѽ�k`D�>P�Ń
vr�z�1al9uN޾�9�v�q�]@3���;��J��af*|�c5B!�Q��QbF2��}��-}��r��%0��n+M�:�}3d� !�R���y�t\8~�8�`��Ҝ`K�/�� .?��B�9�� ۽�-C[w�1@�FO���g�c�����S���.n�5���B�%��gU�=s�ې�LQ0����!�[Q�Wl�ƍB)
pB!�	Q�B!N��BqB��B�� '�PK��ʯ��c�.��_/w�ƾ��sz?B8!�@��u�zL�?G���*�K=G��߀�(�	!�'DNH5���)H�ʹz���D��w]:7R�[=���O�à '������V؋ �!΁-,���@��]�pg�;=	�e&!����Ӯ�0�������Xd�!#�V�.D `$��rFb��	#���3Gٚ<����n��B��������H��R'�R6��bU'�`����[������~�x�O��u=����ͼ<��6ĩ6�B��Q�B!N��4z$*��f��E�U��=!�Rx$ܺ ���w;���}�BHE17��_d?�@P���쿖i��t�$�ɘj2	L2��ӛ���3L��@!�9����d�6Im4�
&6��>b���H,�*b2$���u�Z�1��$l���;��7nDM�afCFҎTN�����N��UG$����G�� ᾼa�k�es�HUuՠ�<!��cb���ν��Q�i%��ai$��+��u� S~�H��ץc���'�?�wb�����T��2�;�6����c�r�Z�+��������񬌩��~f�H���������Wګ<�vQ��B2�:É��I�ŭ��͍!�������A�uPx,V
����Ժ�2��������3�~x���7�>�T��R��/*M������0�O[�9*n�nvPB{��oF*B!���tͩ��α��N����yqKu3����#�K�[���C��m�,�s��~�Oz��}�]g��"�I�`$�^a��F�ɜ��ب�6�w��yq�D�C�tUy��1T�N!��r���܁q�cm�|1����z�zm�
D��Q�^g8����Rx#�W��>�9s�g�]�������fm��=�ikԶ��������<B!�t6/cC\���}|LԶ-sF�zR�>���u27sɁ�;�X;��b��i�>�jm�L�ǋ�0��Y�+z��bח��4#=�R���B��R�Z��뤊��0kl�2���w�y9[Ą�v�-����Z�.6�G����&�\���'>�;u�9��� �
�BH�R����I]���ܓ�`γ����|��D�z`��R����c�<^<M��g�pV�N���BN!��2L��|�+U���~�%�3��նgS�?!M�o2yc��8<у�(B!�3y��P���ypn�>��x[:�������%�da�#�׀'j�� �B�A��~x�3	x�6��h��|�Ɩcm
���^2)����/��8�L���5�B)+�½������L�8f�H߱!�m
�Z�}y��El�e����\�H�$B!� � f?n2���<�T�O���]�m�)��E���F<���˹D�hp0r�������. 
!9;���v�}��BH�sJư_V�q.OF�KG��%���'�}%���� ��M��T�_�gW�<���:bY'p #�=˞��n�f�cx�m,?�B�V�T��$:2Z[���� ���j2� [�+5�Cg�[G"WOpiP���z�fHE�#3Vz1��}B�!�z�,X��.w�ϟ�ʖ�=aNܷ@!��x�%�6�k�f�j�}��nr7�٪#��<;3(�q�֎����i�p	�*]��M�ɖ��y|Ќ���r�1� �y���M+�j��%����������f;��	]?�y�k�Ʒ���>}�$=|����4�5����`�Z���y ��Ok����C�r�����V���u*�fg���ka��N���� ��J�q/F��ҝr�H��Uc��	')�c���4{B����K���k=C@!�q�5z�����=�t�v"�վ/,n*W

�����Q�;�����[��I�Ξ�x؆����8!v�Y�t۫i�=j�Ų<68lp��
�V�P���Z���i!�%dLj��'q��1�=�2���e��T&;�K�]���A��2��<fDx�vJ�Zw;-�V^A�{ܞ��<�x��"�u=l8�n�އ�)_s>�eW	�`0�BHթ)��:E�a�/n^�#�`DX�O��~�����4�)]d�uqؠ���;K��*�!Q/�����k��zH��/�2�����
���yW���օqf{w�:�#���B�X �����LM|�p�/<�	?�c���W������-��R*��5���D��!�RN��wo7��>|���<ʹ-�b��;.dְQ�ŲEM����J�#,H�}w5�r8�~���k����c�,xi#4(��&�pHxYt�f��d�z��K�yc�Im�ZoJ��$
����#q�Ǹ�b�/v�/��ڼ��c0�QMWO
pBqX�\�҄�����Ka�Hc4��I �1/��ߣ
j��@��գ{��wf�����.���LC�`8�(8@��#a�- � N�E�,���]�"k���
n�ʕ@!��`3/��eo�!d��u]T8*�nՖ�D�����۳��	x�H!�1AN!�8!
pB!�	Q��w-�۬��cZ��/�X�!��f�z�߯��ƗB!�(�y4��@n�՜A/�t������BH>f�Q_��Dx�zrbo �B���$nsz��xH��U�	�T'����s+�v�$wۘ����T��+.���C���.!�XB^A'n_�k��<~�?�6^Uh�]B���BqB��B�� '�B�8!��(�	!�'DN!�8!
pB!�	Q�B!N��BqB��B�� '�B�8!��(�	!�'DN!�8!
pB!�	Q�B!N��T9/�+(�2x�djr C��˹\�
�=�Z=&]��!�8�RFot	�Qm����W�2��{��W0���>�;�B`\��V����S8p�B�
pR�$"֌|:�i��Z��0��ТF ��k�L& �[P��J7�Ɂ�����]=	�^>^�ǋ���I�z �T�҅���$|_���)p��z���
�R�P��JW��HIu=|�BlEN*#)���B�8!�℘��JC�{w������5 U��D�.�s�b^6h+0ԆB�D"Bs�
˔�/���X
6#������Xd����i#q�W�R�o�#��r�q���'r2`oF$�@!�TT6	��yC{�Ȅ�ۓa�;����\<���e�������9!��r���ġ�5�����ZN�����͖�[�]`U�m��U!�b� �&֨ތ��Sx>o���k +݁yY@!����\��pm��̩IBx�F |��&\�iaB!�vP�T�.�NXg^s�d�M&?%x���2zC�N��6�SL F�P�Ö���Eb���x���Zx��Vb�V���|���~��`4w���~�8���	�v��d!����K`2[�%���:}�^��g4$�GeBƫ#�qe�*���J�������\�M��O��<��sԼ��|��9Ĳ��uu�/�&��]u�-�q�-����B�PK,��T��'�С_)�8�Z���PY�A�ɕЫqۂ��ܽRp[.��WR'n�!�C�����ob���[���f�x��\�5KL���rn$j4�6/������&d��-W|�X��UY�xjgg&�H|yr�����)��<{],�%������⵾�X&���6�ǳ������d�-Q�?�_~	:�I�Ƿn���o��L	���p$����T79r7h���r�i7�BW]T��@���?]�7��N{e�¸�����
�qk؛kF�{�����Hl׆�Z�n_֣�~������VM����L��K���}6@*���E�굺���=�Fm;b�c�Dm[m�6�D[7�#>b���1��j����]�1�ܽk�g����M{Tp;1#�Ⱦ�H�� B!�#b������H�հy�q��mgm=禅���f;�A���H�ҟ�&7�@Zf`�g{���o�I�,�sU9c@7�O��x��P����1l�|��cOC����T�^�HT��8Z+\�t��ی3�9p��I���:��}���T�P��V�����<�ڰ��i�)2�`0��M�-j���/v~쟢�!��\|�Ȅ��$O��	�]>�q��1V��-�}�}f�ҧ\�������dnc�;��������:;��*����wT�WJ��(v\<�m���:*=,�;���}L����{K����#vvP����\|`�3֎)�ؿyA��&�/�Z[*W�񢰧�F6���-ry��^��#)�N�T�!*��B�����&�+Y��i�+}��,��L�>���w�y9[�Ǆ�v�-���D�f�#yx]pK�{n�G�.�G~�n<{�1/��[�}8媿D�oBy|�K��|!���������c�c�Ŧ�E��d\� u� ��@mjxO�W�_x	�4�n3�$U���~�fn��XBN!�������a#_ϓ��n9���z�*[��)��IS�L��ǘ�<� x��-6����~�9B!�Y���5ix�8�։N�q�Ǥw���V��)�"#��K40��e'�u��^�v��>����%�Rqb+Y�Lϱ�!ee`��lS��i�wkl9֦ oI�\�始�@dh�~��ǹ二F 7_=��eF	!䱧��Z�{#��i>�Gl45��<2�H���wlq��f��{#7�L;��n>�%42-��2�B��-�`����: O.��ql�>��c߮��kS�����'�B1v�[�ǹ<��і�=��TA!�{h%����J>��C$<q�^���D�� ��RY��]wGn��P�^�duc's��F#$R�B�c/Q�-�	�����;�F�J�#�+4�3-@´��I$Cl9�� vf����
x����d}��^���1d��{�]l�:&�ąBwz6.���J�Zb��X"�hr�ao�T���5h6��d�-3Z["w	�9<2z��k�Y��A-�.3�g��nÆ�>x낭;�����!��s����8-�Q.�J7x�K��c.%݁�ΔZ�C!��	��Q��˚�.nQܡ�;x��a�.6��˂��Y�Ӄ~����K�����P;P�:�)��x�\(�U����w�Y��Lc��C[�VJw�[���up���Ag�"h�� �ܼ@(£�48w�*h����\e
Ӷ��c\;ENq*g�LH3谝��>��>�r��C��EE�i��!aC:���E�	��E�J�񌙃�Y�㞹c�x�C��T�o�K�/��ǋc$�N.^�Da�ol^�-�	�5ll{�|��Hl��cW��*�>���s�c;7y�V�\������������BH��j��iI𼷿���b���RxF<asT�[�:k�������M:R_�p�
���3��}��5�E�0$jl��:Cd���X��E	�"�����׵?~W�	c��Gs���%��\�j( ˯�&��AUh�[���<k�ݯ��`t��08�+}5~����^)�B�pz����s !�	���]�BV=���~wF��q����Q����ʘ��B�PG&�j,QTBL������3C�L��(���ÿ��c����j���^�R`�2�y�4Q���v�^\���<�3���e���X\��̊c���.�TE�[&����Qû0w�D�� � I���Hp�w/X?H�	��lL�kٌ�o�͸f��"[Pl�T[���K���1�&�\(��a�51�+��s3��u������޻sj�dh����=��H�{�{y��n�ٛ���8�Y��bR���yL��үA��]?_�o����h2B� ��5�����u��w�~f���r@!��z-�xt��L)�gO�T�nu؛u�A�F�JYG	m�o�:��8e��Gw�b^v��l�η��n��G`0������¦��a��Wa���� '���uY�+��D��N�f�S8^Max߮�eC����u�s��r��	���ĭ�m�p��u<|����KOB!��|n&|v�&L�Q��R[h�S���{V
lKyFT%6������Q��X������3�`F�����+@
pB�|����x��}���X� �*�q:���7#������U�,�}#%���'�����	�!�� NM��l�����S�:U���8��j�Ě��A�..�����l�8�2��B�/}���#e*��?!���@�}�]�NBs�4�*�_"/�dl�[�^՘5Ƣ�n��f����!���.�u*'��N�.��z|o�Ö�	!�b8�t��cVIU%�����!���G3��o�e����o��g÷��J=o��Q�03��;鏠����ng<B�8�pJU�l���AY�a܊f�!�`�=��z���W+�<1���	���B�8)�����|��|��ϳ:a'�n���7��®KǀBlE^A�R����U8M�=���~Y�t#{��̖z��	�Y{�WX�^Ԙ�h\B�s� ��d�x���n�=��WN�zL�������i`�������G�b�����6h!%'����B�����$�����R�{�?Ȫ>�!��P�B!N��BqB��B�� '�B�8!��(�	!�'DN!�8!
pB!�	Q�B!N��BqB��B�� '�B�8!��(�	!�'DN!�8!
pB!�	Q�B!N��BqB�h����{w��A�� �$j�pY��٠5�B�T ��
4���_"OF�bYU� ݌FS��)�%0�bwU|��h"SBoW/И�p"'��'�#�!����K���7�W�q!��É��U����{V
lKyFB!e%g�A���Ճ-�:Hɵ�*��	���["o�p�Տ��mmB!��+Q��u����r� ���Hཚ�aU�m�;/!��Ҵ��p�-q��r�8u�#�P�jԅ�݂��B��>U�� F�|U��1�M�=b��O�F^B��*�t�ސ��<�3�@h2Ʌ���H\Ã[���_�D�:�0�*��u@!�����l�4�N�bбy�O�@ 	k�07F\e��M�w�ss�5�k:0%2K�����9�	C�A;��X�Q\IW'&�uΝ;��Y�L�ƥ�Pb�XȬa�j�d�*�,u4�������u�U�E��Z�>p��- �R�0;����:�Y�y1/��=Mn�օq���GD�pv���2��RU��*���P;��~4�����k�ؕ�����ng�l�6���O��l�)�ڵu?ˠ7&d���ia�W���m��3���!�ۻ��r1f�
���_�iP�|Tp!�g8q�"��=�?��t4�B�B7�3�>���t��/�y�c"�f�w���F�{����g*!c׆��Z�n_v�}�{S�}f���X��/�w'��p=WO���W@�N�;���#n�Σ�>fˢ-�t�CO�S��!�H�3н�I�#�Y������`Q��ˉ}��@4�O��B*��-*�w�����V�I��yrǒ��sST�rmؠcT^�{2�vojrs�e&|�����ۖ>�q]9mP7W�8���:��h:��5"n���o[Զ����U�}J��D	h�p�S9P�4z-�jՠ�ȸ���.0�{0��m�r��}+l=Zj�'��j�p6d���1�g����X����·P�̡�=T�[eB!��:��Tnng�bK�X��x����>���=��v67#nˢ�m�}|\Ԗn�B6vv�cn�[����$�1�{�x�g��ӄ�_�^	�iҞ��r� ��>X��g��� �¿NJw���fg~�=���Y�-�}��l�������E��S�0����"_x��T���Ee�u��"��=�m���z�(/3UMe*� �P����Xq8�۰*}R�`x�CPI��~ſ�r���v��3�3�BH�a��&l&����j5bfRE�#-S76C�Ov��?���h�7G��,�8[Ɓ���]l����u�-���dV�<�ߩ�	=�x���dB!ԒH�7A�;�M޸�o^^�T��5l�m3Saݑ\Ƿ����BH���e�|!�������I[��]��7g��@�[��}�z�-��4�K�θ���K��u��'i:�F�Kws�j�+��V*�u������gF��K'� �Ry�j^��o��{�s}n�<�������W���JW��dP��\߆[��!��)�����@,���.�?�Fw���F$��w.��?�q#5L&7�����{p���~F
����.� �FH�*�$]�����t��/�x�F�ʖ�l
�v�ԃ&�'�1�Mk2� ����Np."ǟd.�T���/�4�6�s��!�mց��g$sp_�o�n����_>7��6{M7����`p`��.X�!	�����.&��������лI{�X���ܹ���9���j]�/����7��3���1�o�$¡+��ʣ;�j?x����E�3{6n�m�{1�O4���w��-x��%���1 �V*��Zm�����Z'�%�p U�<�![:�ٔr����%�d�������Ҋ\,��r�9n3�p���V�`�K����E>��Cq��	l�|�?�>��=\M��|j�z��N�]@Sh�S�Թ`d�մ�Ӕ+][�%r�,��.,9�fΰ6=����]ka�q\�
��M2�,�}�����&~?s�8�iH^�ă�<��`��ٵA���M}���>�.���Bx+�>W2�f/�hD1Gl%Yټ����W�8��d0M[�ۦICl
����ʥZ~��D���|�K��hr��}lI��?�/u
/wu=kZ<Nʈ���;�������F<6Z�7�CS��:V�����ᣡ���cA�������}?:��}c:�iό.�)Bٚ<n~De�Z	{����M��ob� ���5p�Z����Z�{#��i>�G`4�"���H߱!�m
�I��܁0��o7�����e9x�1~hٙ�6�*Y���~�ɰ�p��r�>��m�4�E�_<7�?��3��������Zۣ�*��F#<��I��7���?��5?ު����w����jX�W\�;��`�K�ܦW�}�
7�i���-k� ���~<������uz^6$g���W���y��'�`����: O.���u�J��x�J;֦ w3�'�B1v�[�ǹ<��і�=t�vF,�q�m��P���!��R|sh��ՄXEy�����;�C����� /?�1 �}�vi>a0H	tiЊk�0�܋�n�~�/wf�*�	{q���w�Όa[�G�%�]o.�����|X���A���&��g6��l���ݫp�-Q�z��.\eJ��l�ZdD�X)U<G�\��/��	�%������G O<�e�+���m�X6�+��1�uw��
%�1N 6v2�O�^}':��6~@hх�q>�U�X�9�����l�ݶx�o� !l�~�ʿ�a){˫�	r�ah�0��)0bE��ϵ�cu2����k$��w��yA���F�]_xpe�A��mK}>��gK�㾁��%�m�/.sxc���7��:a��կ��17\��?s�I�0�^>�����J���o,�P	?v�{�O(��
F���] ��D�4�ߖ�L�X]��shD�$:2�B%�a�s�)[O��M�[j���5l_�� \��W����\���Vz�=��?{I�]哸 �p�/mc��G�ׇ6��	�ټ�	��~�x�p/���y;�`SB}/��Cr���нQ�Gp`/�W6,�Jҁ��S��\|~�i�o|
���f����Wlֈ�24�Y���;<��ۿ,�E���|���ǝ�I� ��uز|��Tnź|�{-��z���ܖ����'\�`��?�'j7[`�o68y�<�z6|?�Â��o�ퟗ��?b����a-����1���������V���Nj'�\��7��b�:*�u�5�
;0nc	��}����������, ���q9/�4�y1�47{{s|E���U�=_�� 6s]Bg�� v���x����l%w{x�Z�2c���N��'P�j���Xv:T5��(m�Տ	{������`��	���=0������X|�v��B߃'�熁!���X�~�;q=˻4��jI���'�w���b������EY����'�O���lI�_X�����i��SJ�̈́���������N��a��/�y�=ȗ�x�`������7����.��0m��\`3����Ě���͑�R���!b�
H*�o��O-.l���6�矣p��i����#3Vq=��
?����}���6��3�{��y����XN�� G�U�c�Ç�-�t��3����VK]���9����������f	h�P�����8�{[��fmؐn�n?^���:�U[�b���LP
���\Mc	�x�)�6Vbɡ"�\�`z|&��R+V����S`ǹ?��0�%v,U����:�k��4��b�	>ǨU���a@c��6o�Z��5�9���,q�(����/�r��`?�i��U�����d��\m��?��"���������u��n�5�!��O�"��|�T�	�V?��7��^G�S6-����Tp�l0c���W��º0l6�?{�Ś',e{M��Ռ��j��E��{�c����H�Hb�Ss���/�,u�ßkP>	y�k����T"�fΰG�z��M�BF�F���n��'w,�Z�M��uj/w��{!�)��Z*ǒ����ǻ͎6ཧ�]����D�_�ċ����x���v�|�z���V�ҝ�\U�3��,%�U~�gq��a�4�JL[�Rn�:W��FX�U�8��9X*���	nF<k3�e�W���R/g��[�����eoÉ��@)��������q�j�x��"㩋æ�^~v��R_�5j��̂�]l/@����"��+=�ߋ�7^��eP���r�%�5Y
ot��e������-�c��Y6��]�`�莋l����V��ɵ���3a7{Q��W-��kH�Ү��S����7/���.Ue�^O*WI���d3��<�h{��"����k�6�:��_P��"b��T�_�G<7�V=��$�L/jxXPhm�|aS��� ,��k�q&������
澒�{�����X��཯��gs!��y
�ʆ%=,��p�,��Î^ϭ�͖�Ym"��m�/�J���d��Y6O����|����)M��\�n�]"�����p�5�[&/�����*p�M�[����]TP_�0��]$f��{��xn�=Cn��yq%&ڈ� �9���uĲ���ڕ��'�JB�k�5�5��#O�����}̴�/���J`j�)*`��
�7��\Y�ݾO7����5��&c��
R��È}=I���r٫�u�w�A
�\i�Ɲ�KO�k5����#;�q��a{&��ƶZlS�T
�J�ۆ�ŝ�f�~�u�BX����������-sV+[�)��Iep�t��U�y�p-�Q��|\<`�?q=�]�J�bHPbW�s4�]�=��aGF
��?�%݅0�w+������ʆ�A�~�X}�^�@m0��<�c�H�����Y�4X�~�ŽK�fn���	�I����{L}�/�����\��Pz��k��ې����#�Xj�
�N�Dk���ɢ=�s�ٱj?��!��o�~Qb�Ql^���D�揃Ӻ������V�̲��m��\���C���]9�<��@��cp�����[�Rj[G>�\�@�o٬xӷ�̨5Xpd7���/0j+U��Jnє6���G)�F#�J��胅�vP�1�Xn��!or���4I7)����wm�*~�f��㇧��:]9����-S�b�9V�[���f�>��o�aV*���zz�,�.5����+�TOWجXɆ��u�j�s�:��uZX�|�h�����w�8WҴ�&����|�N0�{/}�`h^��j*�����8r�m�~|��W�0��c¹^��`���og����x�懦>[0|�:�eMͭ<��8֟T_��`��w�ۭ���9e�M ��R`[�CP�h}���ׇ�Xp4��nӹ{�-0��2��qY�u���?\
Ǔ[�äp6@Kp��CWN��:�7���>sp�^����@*�6�wu�u�=\�@X���e�T����΀��I��&[x�`8�����R�8���#;��N��څ��o,��c�a/n�ñ�,��g�{��u�8�^��VX�?���Ǖg4�/��!>+�q�v8��U�3�b=w&�^o29D������rs�^Vg�v������6��^���m�pSt�8�:z��O�[��E�����'��J�����Y��$78��������,�~8Do��y<<�i`C�=.�[�U�D�����E.t�@g_��h,����b���f����q#�>U0ovi��z���*������<�j�>�!Ǫ���>)r?65D�X]��s����(��z/zi�,q�k^�2�/xp&;kp9
��O�dr����������8R��M�5O�mfu?�ȅ}��T�
V�NzYa���c	;�m;��]�����U��j#�І�Lݼ��)}_0���6?�Τ�O-���+녇�}�����/�pQ�w�]�tk؆k'�c�ZB��N:�m�-��H�y�,�AKʧ�[pe6��,�����g�7K����A�u���q��8�<�o]�Zt,�>��=�l��{��[�65K�����Qf@�kpmp�������f	v���b&���Zr�VyB���Ɉv}�5�N�A����W�Z��ln�H#������P�۟_�t��c�n�G�Ꭿi��EV��Y�6X�[��98W�-cǫ
6mlٕ[����[�������A�~ŝO�N�o��(���X�3�0E�o[*^���*`4$�;7���Q��8����-ځ��-�&�����������>�*�/���"��u���=�[y�zpD��:.؂�EǕ�6���kM���C���/�ݷ�H��ՏTO�vr?���r�0t �*����gk��Kl8{��',���=�I��\����-�c����8egU�չ��K�iV{5iǍ����I�u�[��Q`u���n�F�зYx��ƍi�eV�.�8���J/ܾ�/['HB����u���ʶ�o萋h8��v���ힲ8v7.����Ϯ�����{/�v�qKo���5�Ly�ynyͥ�~��*�$�;a�Ҙ֎wX�?��x���\�4�8f�ε���Z*�\����aq�Όc�}X�R��8
p;�s,�a��������|�T���XR��ޗ�s�d� ��װ���ۦ�ӟ�-6��`��ލ���U�),��!��\p�������_�0�1�1�1�1<W����+�6����s�-�ʲD'NG?�v4a�\�c�Jn�V��ߵH��$��̐�=�q5.졌��o�<���ζ�4�XJ�iGW��OF��?�z6n�m'o_��v��FTf�㒣G����ڔz��W�,�pV����sO>S���n`�A{�A���p�S�'e$�{p�[�g���]��8:
p;�޽���'Dr�m��������WN�-X�+w����X�����L0G���om�壦r��8�-�Տ���h�n�ze�ћ���o���������C�p��)��UJ�o�k�ㆰ�̬%�s���O��� ��:�pp�W���Rv���a�������|�2w��?�z���%؉K�8̨��~�4�ث=B��q����M`��p�-��|�M�bo�������PY0�?:	�v/�ЉM"�~�>��}��7��U�J�ّ�_�8
p;��޵���҇��IsD��4Wx����a��f��QU�8����b����׹
,�]o~�]<�7/�J��bk�qe\┥s���i@�Ifp���l��V�/����O�m�&%��r��]8�8
p�4p,pP��ő%����[l�*`[4.&���.���0hV�.w?־�����='n���*
��g�^pb��/��}F���Z�8����>�mgCU����^_��2��5Pt�,(��?��|x�U�Wֲvp��;���5���5ݼ��ժ�&{�?1�aǰc�?�Dqӳ��r��,�oNn��%R��SI�7l*�)[?�
x*]��&#�#�]/JӤF �|s)��m��yp3�,(��;�\O��_8�)~O��|����?��\U0�qX�ܶbL8t�o�6.��Ӵ��П-�~�.�Sm�t��8Kˊ�דu�sV��.<s��Mxe����Y�J��0��n��.��Y�������8�1�X��gK�U	�/�X<��}���&��3^� ����د��a]�{�ۢC�� �Pa�l���sDAgM�A�x�F�ك����
?N�k1��ׇ6sC	q&������iu?./�m�Xu~/=��qjx���������tt��08�+L�^k�*�<�O7�`�q�@V�W��Ҷ7|1j�+�c�qli��/��a�}ӈg���'�bj���V��"��B�8q:��N�1?�U��C����:-z	"�N�fs�/���֦'L�U��8�Mƀ�.0�]�j���D���)f�#�pl7���b���G����13��΃J�������� 'N��
U�ε%�w��Hc���*\s�5�m���s~x�#n��|�8����I`l�mꥭ�^�ܡ�a���2�P�$1��EpK���EǏ���#RHd��Ԫ�����\B�8q:~ؙm�3����i�T�¨U�m^Uٰ��݂�9�Ϡ�%䭯.����yI�3��|�X�]���4�]��\�z�����-�֍.=�#����N�=it����~;���1 ��P��4g۷����GG�&|r�w��Y�tfa8k���sC�pu����N�2��<��0�G�9X����	l��^#��ǖ����1�ƽiRTA�°�`ܺ��tx�5�7�aB$7/�%8JA��*t�|(��SR�\�o߻_@m�V���~��-|�g�ߵ�!'�����m�Nݹk��.2el���X�Zxy�|�9�"�����D��,>}�y�q��_w/6O^Xb�v���w���q��`SB���0{���
���B�<� q��i]~t�/�Ć��'�ȇU����'�����p8Ybz2lyu!ש-�,���yХ~ L߲Z�jKF��
��U8f�p���S�N�_>7�`�[>l3�f�;�U����a_	�V��ǯ��m��؂�85�����\ ��s����%��7�~-��'�9p�t�d2�|�S����w��M'�C���a�==Q0�+�pL�1��1�#W�ÞG�����/nCM}�r�	�&#_jn&�7qz����Z����{^ٸ���_B���CX�%�¡�ߔ��=���?ի9i�Y�wٛ6�x�p�ql�/��Q� �"(����ad��@�H�U��TC�㷋���!/[܏�Ͱ�yp�n�*X8�`��S���S��Z�>U�Z��ڀ��8Mx3B������^�w��I ��Q��I�杸�=h=��]�u�<$ܺ��wm��Na`�.\��wGvp�::����7�x�Z����	���������_>?�[�����4��8;ft���J��z��!�Ic2B�N��<��΅yY�6:�bj������D ���l����\O���W��r��cgqs�ώ��刽��ү�Rde�w)_=�.�VC��m���qsw�����!�ɄBh!s��2%�K���~�Hy�kR^��f4��2R=J `$��*
��H̾�
���Z6�O�f�o��@��k�&�'ܖ0T�aoX���8�RCa����R�د�fG��
�(�M��Su�w�Z���I�|�gJ�؇��?ڹ)�O,��n>�N�
	l3�ÉH��.*�̖������o����Icu��a���p)E����"+݀�>��m���n��)RoS�w�w+_)���&M�����ڑi�����<a�)��+�J6�j-$Ϲ��q�˖���^H
�;�)���R�b�g���j�H:��&Y�}k�N�׀�9���F��`c��C�l��Y4��&�pq����G�.\/dd%��	�T OotMO*��BK_?�G�H�6�nu��%6�3�N{Zwv/q�a�s��U&M��z��K��[�}��W��<��#<yuZ�z�X�b���6�5�A2u��:Ѭ�|Ƙ�����H^�}�)7y&�9�%l2�'�Ax�g�˂���0�6z
��>+�r��,�X?��d����h�����ϛ�
���W��%�m����,X�"�k�@���Zmh΁���@�>�S�|�����N"%]�W�\���^֝�� ��3���?��ea�,���>���$�]Ëe�smd#,���Y��gz�����m�ގ}]�y`�h���3���d (��9�3��dr�~�|�Z��uw�𵰰h�w���5�9I)b�L��୰����]
mBvG������1-��qobc^Gk�Kg���3dP��x*Tk� �˜��_ܣ�������e�'��U�<4���&?V��͙c�4���Č5�Aj
g8���|� �O?��z�t���4�YJ5��9�{��ʥ"6��ԡ6e�2�v��������$�Q�>q��]�&�m��Ut|�[aEM�2�L�����re�%�Zῧ�c��i�)f�,��n��K��9�����*������NT��'��>[���:�{\˶���ut.�����NN=2�Y/��ù���̧i���^#ta������u�$�%����oF0rk��̣z��[4�grv��f��O
�]�<]��,�=3�b�B�7##�>���m��s�����^=���9���x�6�����:����e'>j ���:~�n����þn]�=�lJ��y�T�p.,���)��ubZG7��յ���2}+��jG֡~2<m���1}�j6�4�� rR;��_p����dl) ����D�YZ3ų�ӣ�Q��c���%�z��B@հ+4�4xY�|a��<��k���ظ�!��%��l�X-|Y�v��\�w�+̚�>�Dk����Ԍ�[�ߦ3��oK��FE:x^�k��d��6N{&�}��S��^"o��*f���
nN�2��j]�4q�Lg">P|�s<|��<�5��B��s��VXxt+�v�����zVk��˗.�����vR���6�n{�m�+���L��ǆ/�	�Ӭ��,Ҝ�׹���B8M���Ɂ�9�>��]E����1?(�76 G�*.&�RDL� �@�r���Ώ��le'��J�YZ��DD�ӄ�8c��9d����S�~�i�WUW�⢧R�����#ýM	މ옹��ҧy�j�����
�L/��J"C(-A�+�8�����h�_��j��YC��LAt�w�o��x��5�����Eh0����BpJ/C�2�3S�|5��P�7f�j��f�Q��͘��gjF%ѫ��ك<]�]8��f�|�Q��Y�z�R:�(��|�j����NrJ;�2Q0]D$�%\
m45�d�`�0�(�6�ݔ��vv����j�χ~�tq�n�""7��M��:�Ռ����|aW�B�N޺#����~�y���Ξ]u�^��-�8�:A��N�C���h�B��+�K
��ן�'���]�ΕQǊ)��u���u����J�M���1���BV�0���GhӅ��裒���ˑa+��}$���ej�6�qm�WrvkAr)"lꁙ�.*���l��Sد�\jiJ�!q������qb�^���o2*?�P/l�Lr�����l�����m��b�b ����7�����eZ 0ـb���#Ȓm?�f��I���dY�?/�����X<�\MzN��Cۜ����	�b�F#��M�s������ǽs�+$�V?�D�o�0��yb��ڗ�1;� �N��E�b����eChjg��F���v�� ����+�M�.���ꏑ���禂���S;��ZƌQ`_��/LG�U�$��+隞@���18��!S{��S��pO���ll?��DR��wz��5�<�[�kћ:Vhht< x���CGٕ�L�[�5Q�6��)ճǻ�ք���ZI'��$/cb��9OT��V�D�"I �+����Xx�����8�"�&w'�f�Q��^&5�a��<�H\B<�z��c�ҽ���b�^�s���T`��g�v��w���q8�ȢT��C�f�T��>>���w�wD�Ҋ�#Zm�b�M�M8O�H8��6�͋�q, �C4���XJݪ4!�R��V��)ڋM+ >�R��;���;l/:΀��*�-Κ��(��vl��7�x����\U;:!��T�+�$�a緬Z}$HĹ��j��GϜ�_k/K}��,A��$B#wѻ��bK8��@����B �K;�f�y�:�1V�����t_h�o�t� ��v��nru�JL��D��uޡM'Nr�b�cX�d%�<A��hm���o����� >df;�F�y�<-��N;Ć${��i���PZ��f u���*X"�@�����(BjR��wGػ��l��m�~���v�9��w�Z2S�#w.�#�X�@��^P�rI��ie��x{�\������o��=`Q���ؚ%j�U&ȱ�[�ǲKP�5��#G�۞���Wk�|�
�I����7�U\Mf#�̥9����M�e���T^/�� 2�Y�Z?��/�!���Wl�j;tZJ�U�rR<�q���et6U�_��Bы$�C��=�D� �����^Y��	�z��Ғ.cȻL�?�ٱ����/�ӍX��]�eme����h�Y��#3;Z��K��2�V�7�N�XLJyL��Mc*kK��eNzb�k|��%�h����h���Ptl�l�C�;�sS�̹L^ �q�Vn�z��9��ޕ���I���ӟȺ�䝅/�x��I����;�*�gS���D�Q;�l���m��y�ھ��s+tf���z�;�9@@Z����b�}�_����O��[gY������ȑ;����?�����g��vZ�f���`���&�tv�xa?uX2�$7��|�%U2��U��E*���b蠐�O޽�~ޱ��st�\X@�1A�c/<�ڡJ;�v��"�������{��d&ٔ��Ŝg4���i5%��A2=t�g�_%|�����aK28x��ƻ%\`�ؑAGW�G��4�89���3��h�f49gݠG�J��\[� ���fs���>�A�a��%t��y��ǟ9��B�P�l�
uT/p,8��e㍋W�>5ZQ��Ռ~F���KS�E>�S�/z݊��R��{ @L�X�6U�b.�ծ
�d��9U����zO�8i�8C��_��*Y���tk#�trm�jL����Sr/��%\;����2�� ��j���B�Q2{��&�Ŵ��ӷ�j���9��ۯc�LN��,4��5M� A�����3�>�u_3��ןӟ�G[h�=�/�<���e����%���4������}Ɓ�ȨF]Y07Vf�[�<����L������BL��AiG׮a>���o9���n�ӼU)'ɪԉ�rp��r�n��z�*�k�����I�RR# ����F7�4e�i2�>-J�qtݡ������+2A�F�q\Ӟ�B�u���G���q�ӶE�Iދ����md�#��N���,TJ 7�K,������dQ��BG�-��ԍ�x�7#���ޒ�_0����P���R������?>'�I��PzK��ϋ��%e�vi}ZT���)��=�E�rB,S�䒏��U^���LȰ��O��)ލ��Ȧ�k�x��jF?pO�JY�5�	�x�!�������ի���7���!o��|�f�e]�Q�*�.�0Ë���o�����ƨ�9���g�7�M
ޘ��|�YAϪ���j��@a�˟�t�^�!� ��}�Ne=Ɂ��d�~��M* ��~�Xj[n?-�4ʠ�v�W�֋- 8�2�����9�n���J������薽7M	�ߘ�����Wtr��,W�Mt$���I�&��Ѥ������I o?�GӬq�?�W�++-0�l������k�	F<�����:h��}�to���)��aR{Ǽ2����
��t�{�P2O�(��w���!�Z�ӏ9R�MR�A�2�,9)cL�lTL,��N}V���)
%�yG��,PT�֞���TnLM�W��6أ�����~I�4'����^�؞�>�4�{��1����|�d����A�պ�$�
y��˲�����͘�S�%?�ח�E������Bj����ȦR��=�m-2����/�>�������'�ܭ���ZYAO��A���bn���s
ǲ��Lм�J�{CZ��An�9�R��]�4�lO+�������ַٿ�w0]@�M�h�T	��'R.W�S�&��^���f��c���Xb�Hʎ���A�6��}kɖ��']��?��2��t��UI�� ~��m���{^�l�hEw_�Z0�,�%���5wy�S�� 9���D����Kޯim���V�"%��J���"��B����²A��&'��.�K9{�h8>{�{M̽���g�|vv��{�i:ԅ#��mVS�'��.~B��g����NTS���$x�!�I��8�������E+��n_��9�����,��:o� ɅǷȖ�6t�u��a�}�3���~��`A��:��eZ��Aÿ�L��J�W��q�#���c�%/�2�+�
��&|�����NN��QR�ߒ�#��B0߷D�@0:fMT�S���+N���vcY�A��t4�#��/�4뽽�x�ق7�lQ�E�����-8���v�k�{Я��-ug8�����D-K��{��-�PЕ�V�W��w�#h��G�+Sn�6���M�7BƽT��h�8+�n\�W�J�V�J>(�(�6�1�	�Th@MKTu.��Дe�����3�]��%�%�E��Ƹ�����ϲu)��Vǥ�����T1O1���:uf�#'��B�7���.s.ʨ������dd@����w���+�N�NӒD�j��a|,�Dmv����S2v��|
���z�u.\�z���,k���L��F�������fKdq�4zο�i�f�!�� ~y�jr�3���ӥ����>�5Q���.���J���c;+�F6�
���#Bho��}[3���UWC	�hּLi*)�J�sI��;>c
p���)��b���$�A6!�DټT����3�Agֹ�`#Nz�8��r�'{����t��cI_�ן�q��s&��K;������c ����s:L�2Q9G7蔐���I�-�j��Z�����6^ôloGG�ͨp��	=y����;Vl�Y 7��5[}��7k2Y�1��̋��H� E��a��{���Au�Ӝ�- }My����������t����G�R����a!��]�O���ױZ#,�7�^PQg*l��-� W����M�:�q		��fŚd�������?�C�T�����^�������KO�o�nh�B��Ua��B��ሣU�ڬ�\ȑ:#���m�?Ӡ؈!���{n�#k��i�L�zC��LOv\;.��AEkL�td�����Ӗp�A� ^�e��{�>D����ZJ��L;=���c)�b�����sY���⨆]il��m�e�Oߚޢ΃1	����y����D6B�Rа��̘�Z�J�kz�Q���St����F߯�"�����q���79�Y�H���fd���1�u�:l�fC�It?���U*ǿ]ɹ=��H!h��Y��$��K���@�_���E���h I	dZ1�,V��l�Z��g�]C�-b�]�^$T�J�J���}�;TӠ�/�������]�6�~p#q8���H���j�cA`f��$Y"Ƌt��;���5�8�iU��(�Pt.o�P�v�~�{���v����2��8|I��W����2� ������R��}�Y�����ئl=�9���LTl�Y4��k�i҃
f�i�|\|��@X�cMJT%1l�t�ʤ���}��SA�<;�O�_<qןL���ʜ�-&�����h��`A����b7�>�X4�<��-�tQ-IV�ϝ�Ikx �0Ȁ"[͂��V��,�AY�������e��\������l�f�2���-��2:�7��Jy����φ�u���p~�s��c/�C����(iuA(ɟ��Z/��Yq��������+A�n�%���܂ ;�GZ�g�/��;�����i}�I��,	DIp��a���]�NХ�w�H\j�3a�S:G!�S��-R�-���ݚ�z���:/�)U|מߧ�!z0j�8'=�8']P6�q�3��.��Y���i�wI��RJ�(WK"��|����{��ބ�g�U��T+����;^.�vW'&s�/Cv6���=�Y�㦂&N4��n[L�v/O���G�E��uQ2�xqǚ���.�}�.>I���ѥ]�Q����Z��2hs��� ���z��e��1�l�LMih�,�� ���x�d.�痖�3C�n��Rԯ ;^}\��
�c�� �I��N�lj�̹iK�)�L���~��}���)=z��B��)&VC*5y:�Q�Y�D����D��>�5g�f�d��m��c3b+% ��gF/#��蟗Mz�w^?�{\�n�?�cm� �I ��ᾉ���VkAs�aNa)�EH0m�p��_=F'�_a�)ƀ�z��Y�k�U%�7��ړw���mH�SM���b�Ӈ������\��==jAZ{�o�S��������p8� ��t�W, ��>�:��[�5��f�_G���2Y�A�8�`r�1D��M0���)�rJ�8P��fk�3O�iV���n:��T	�-x �x ��<l�E����;s;g���`ox��ߙT��z��z��L�m�yG|Ҵf.P��	�O3��MQ��=��yt��1��`r�w2z��T/P��/�3:I ��,FM1a�p��96.�b�ӘX�3�����pjY��ɯ�u�{���Z��F8�g�e�e�u3[Y>��,G��%����giC�ɢf���gK��x ��2�>D��=7:N�7��;8�c�� αy�
��sct��c0��7̆4%��0EA�� nN��q�|uO?��+��CHe�dI�>X{V_Z�eu�����X���ъ-��l�C����Y)�1 �d��;��X+<�slS.ƘNs�ݫ6�a_wJ��'��'l_�$N�Uj�ņ��)RC[��"i�~�Ńw"ѱ62�FX��Q�}����_��kl��� )�\M���8��1%����g��ѰjJ�X���ݐ�L���E�}$y��gv�G�PZ�E��M�2S4\�"�k�&b�׹����i&N�-}dtN�_;�cM� αiPN��z���qQG�Tj@��nti�%�R����"=�����7�"ka�ֹ��-��rzR Ŋc�W?���������[��4�� ݲ����U�H�=��KƦy�NdĖߙ�|j�_��Vk�x�U���+��́��3-�4���J�����@�t���s��'�N�c!<��#�d��FN�t�Ҍf�h���a&kZ� ���9����Ƌ���.�6Ѐ�q�x�<n5�G7MKT���GӰM����p��- ��}H8�����y�ѵrf��w��y/��b�����X �?���,(�����tk�Y��Y�bB+�;X�k�ٞ��P���6����<������2�GS�v�����o��f�[G����fg��T8Kn�>���h���d���<�����������5���.��P�R5���2f�}?�Κ�W���
<���v��3a�D��3��o�b��#��w���WY�R�bU�K�Ƭd��?�͏��b�Ń�!�a�0��>��P���GQ�1d�l�r�^��3Ia��P:�q65(Z)E����Ĉ�`�2��[��c� n&P����d�^:D�W�3�����es�}Oر�w��<�w�H�t�$t�8�-vLa��}t��e�VֳZsrH��[�x�5��d��}��s��
t�;��F6�*�>X,C�=����Ol�=������H�r8��f�a��Lh�}��-#j���o��T�py�Ǎ=�]�OҗJA!+�{Я&o�F����v��3�YR�?m[D���'M
������>�N������Y����������$:p�LV�Z�u,�75�j�8y�r�p���D���>~?>h�I�BP�B�8:l!�xD�Ҧ���\��(��P�H
4�o[��A�2��f��2> ����=?�-�@C���?��`����B-1x'���Tzb&C�qC c���!m�x�8k�p3���Y���M�����>�ߙk���>v�l�D���i��`�'m��h �kғم�����lxw�}��M3����dk`+CL Ǵ�>���f�h���PVR�J�vOן?`�p�5���.Yw��#��D	�D�p~����t;:�nD�S��:G^��*����(>���}��K"-�Th �\,v�E���V������s�FF�bo�?�-��,&��yK��͗�脐Y�TEe����+p�{��A�6��l�=�*L�aPW��~p��S1!�*$|�ٕ��Q�"���sQղ ������f�x���.WP{G���I�B@?����+�W��e_�
%ʔ�n�~l��q�B/W�ݣ/��L�H�ƟYS�a��3������@PÛp�:���ug��(��ݮ�߽�2:��Я�����Q�5���sq�/�_�e�rNn�4�U�9�� ���U�=���;{O��_Q���Z#�o�e{�9=2Ӡz�ي�p��[��Kc~Ǒ,��b�78,B���ѻ����5�[�(w]�[�0��_xb8�N�ha|�8���1�{�iS���QH[yd�j.�$#�	܉�T Oot!#/��BK�<��V8ˊ,���Sh�3�_�֬�7��FQ����f6d��_��j��U�׳ =�=oSx��%�2dŉY}KZ�J�X]}�u�M�w^?�B�s���W&=�ƺ��K��Ի����mQ�?�'��O�H�f�I�
����� ���BI���%o�еH����rϕ�!��<�w�����L"5���1C��9А�oݴ4�gN+�<�K��E��2�-[$�h� Be��>�On�(Df'�X�
dc��G���T��ݪ�tt�B����KV�
y��I��S��E޹m�\��� @�L��׏韨0�$��\�10S� ���:ω�Nh{��2�bTXL$�8�>��m��*�x���.�b�loJG���
���Zd6��=�*��ܡNu�0`�?%�9�ͨ.���м5���|ϱ��;�wB�V�x���Z�v�L��A++�A&sJ��}\lܛ���1��o�2��^n��N��S�V��\� �˔��<�G�qK�\6�?fSA�F�0@0��8�l�ԛ�ٰ���P�@�<�@\X<|��l��"�Tsyd&[��^4��S�����N��&�Qf�v�6�$,p�d���ib��k^D�'��i�2�\�!�B��C�L�r�VKO�#�Cb5wb�)f�,k�xc���挋�P@��������߭�ȇ�b�Fo��^�9�}��ʦt����K!;=�;��{A|��19��R��0N��;���4q��imy�7����\$K������V��ħ�9��߅,��f��=�g��4�k��$�=2�"{�-A�b�n?�D���M��M�ѭ:�W�V;�T�IH�k�!'�<{���'�'��'+��1+�_�TѤU]��9T�f�����?��f��ņ�����}�:�wr[�g����.�t"�2#2yh����߉�,�u��l%��7ϦH')�.��SX���f�+�<TuJf/h�[��}��3�׃�iH��z�va�;6p�h��՝=)��A�� _�yJ�A��n_'�\\�ʕf�v�i�5�޽ob���:�����6-����z^���Y	���^�xW5`�т�[������T�)�|�ZgN��t:��[��:�ܳ[�|�o_39�N-�.�p��E0vW���wR�.g���g��Q l�@3�G�f:o�7Am�}����m
������x}!2���)���@� ~t���=OfP��d��D�y[�ܜ=Otݮ��q��G�#[Tv�+/gP(%�9����^�h8}��n
A�oШ��j�yt�S|��AgziW��ed��jJ�������Τ��������T�[�$���%������ֈ7���/�m*+V�����My �-J;���Bw��H�K�������M@*��]��}�����u!ɍ�R��,��܌?8m�uO�i��2�H�®F�N߲3���t�u�������u�^�ٍp�I���rDkUg�~G2[��o\��I�WMЄ��	Cnr.��/���L\��]�"�c[T2�}p%*ly����R��['o��:�uP%g/��+Q��M�ipn�h7�f����~�40��?w�T�!..>�}p��>N�R��m��c��}���ά3=^˛�l�F"�϶+)�;�CA���>�5����ޭJ��/�[�Đ�)V�����݋Ԫtm����U��\���A���Z��N�r51vr���"y%w���M�j�����͓��7v��vx���B o/��ǚ���O��l�ۨq��tg�g�]�vv�]��'"U�8i4ߡ9-��	i��c.��(���I�m����E���eS�sy<����Q�g�! آ/�c�d�\#���s���>��1�'7Nܘ�Q��~kB����j)��I���hQF���B4�ّ$�����D��_#|ѩ���p��G�����@iKY\��KCT���Q�y��W4k^&�p�0�
P�GN����>4�P��A�.Bl��	�}l�f�$�m\��9YQ��"�V����y�!���,^o7���[��
�r"1\}vW��S	&�eX,(�f+Y)��1ޔR0�x�����ē�
�w�<1x{�,��c8��'Q�q�u#���I۠cR^�:*&���GϜ�_k/K}��,A��$B#w��i)!N�)�I��T�]��2�ռ(�̔��f�0������;UlHk��M��j*������pc�k��SI�X?J�a�y5��	�d�		Z??qe}Q|��vj�D-�v����R<�*6�09�6e�h�Ђ� 6����[:�p��B �b�#�ef�i��VߘU_�\� �ɠ�`6}��^Ǻ���*Ѹ��H�,����x{�\������o��=`Q����]�iQi���e�$�� ��ﶰx�m��G"�	.3�2zN��U�#[��פ'e�n<ƴ��}�5���^?���A\ �]�/C�@��+�t������+�w���k�\Q܍TߑDx*m�/�x,w�����^٠�󗊻��	E�<�����Lu&gwɲ~sP8sn�Q�{VJ�]Ë�]=*٨��`�ei�>�0 ��[	�U
��Z*�Y��8f�U��D��N���R<��R՚$�]�b�$\�]�Ny�L2r�;�����=���T]k�v�ϣ����hm=��6C��j�Z!�E�x��F��Ż{�f4c��Fе����d�I"K������4I+Pm3��&ģwS�T�4�~�3�6�sM�1A�c/<�ʾ2b�a�jC4�m�Ge_�$"�ʾ��h o��55��A2=t7�B��\)|�25��;6t����Ϋ���pJ��d6CxL����.ų�`h��4��&���!k÷y/����䏋�CP�TkV_���X�][�����@Km G������зı �u+*�J��ɨT)sG���V��<G��UR���T�;�����C��G5+]��m(I��F6�E�.c&��ӢA)'W��ó��[�D�0�����݇�p����?��E���D�:O�%4�I
�+�iguz��֡1����(�����j�h�$���3˻�Ĕ�Ā�Mj��f�fPW�p��l���tt����<�?p?� �q-ۖtt��J�H)'���5[�w���z�"j�m����儇�F& ���<6Ə��8)��)���U����vG�B�_Wp���DX_y�J�,�*]���Hu"�	�|����E�D�ٜ���-}�s0��÷�w���z�����y�Ѫ��IA�R5hc���~�X�ĥ��˄�M�6T�_*�ω n���^�v�Jo���:����rYG�4ܫJ��@�J7^c����w[���%w�boY�S�Q�J���C]����F7nWC�&���l�
�����Q�h�a���s��c��/��:ex}����ڪ��y���P�U������޹R#6���x��a�U�o���q� �2dg{ө	(p=3|&˺�c��i]����s$�J0�����7�:,G!Q�V?Nݫ43�ڀ��6 ��ix"��C۳a��A}���I2+U���n�c��n��D�c���V��}�.WL��c�褖�oiG6�xd����J����=Zd���_����I���g�Ү�[��9't�T��F�a�a�ß��|}��j�W�\r����szYw�#�L����q����]N
�|o�|�J� e�"Y�|4�@�GGp��9��ܡ�>�_{.NK���rIUu�j>��L���j;�m�IiE��%iǀY�DÒ�d���%������w�Ԙw�1�bp~��S%[��~E��!��I�r,�)aAW�Ń��q"�I����O�0�YL̸���~~��ym�ڊ�����&T;f���ΪT�Z{d����6g.<{9�����oS���GN���D��e2�J�A�Y��9�p,�w[X~B�7Q	ڷ��&��U
U��
�/*BȎV?#kR�����O����鷃�Ľ���L\ %�jJҠ��]�����.O��1|�o���GX���Sng|!�kJ8 U�Qt`�v�LX�Oݳ�,M�*MiQg�;�ł���>+h��_Ye�ܒ���v��^�Lމ4)Q5����TjN��r����(]��	��^��L3�׭��s�X�!���!4o��ゅ��d2)ՙ\���T
/���{�RE܃��+�Fs?..�"�̮Y	��8I��&+\P�~L��g�;���X�_��^�/��֞�/U��~��evt�x�V���5� �O�{��y6�Bt��.=�mP�:�E+����)�TX�N������o[h�p���2�T�`����'tW�P=}��"51��êA���YA�Vi�_ M��h[��8G�����qpy��԰h�T=N��S�g������=��&�m�}�E�Q�,�XP4��B!t�J#�'x�9��M!�m���}�_=f�sk�y�gVg�[k0x'��Y�F
Y.��KV��'wPz�!bx�"�XGJ��񙤖�Mz0��+~�|��s"`Ӊ��p�ͳx��	�#A6_9_	����ƚ�Ā�zy�jZvbM۳��yFR��,V1�m(x�r�er��OLWm�\����b� ���>��.w�#Y�)�^�Q[���k!s[��1=�Bі��)i�}����;P �м���P���B�s�/��Y��,U��a�~c�"R��xJ����߾��m���v��:�@t��Ev��X�� \ӷ�7etv7x_,L��h�3�p������c�
��$�_����6�i]�������c��cf]�q,Í�p���>}�97eRخ,�Mpt�yG;C^�������3(�bk*��}[�$D�\hQ�c��2�W�	�=�����<�7��$��B&��v]?)*��%��T��u�&ū��E��������~~c�}��-�ɻ�3�X�b����.S��R���:v�2�~p�=�����P]*��+jZ�sS����G�f4a�b�ާ���2{V}�:-���
x"$~S�ߥ��Y���'ّ���Ʀ8$R�	��!�l�ۚI��T)�e� ����X�)���ʥ'�ȷ��,^�h���Q������E� ��Y��#c�n�r��hX�2�2ŬF�)Q*�߽��J�c�;���qM{����D5���q�@� ٪&>�i�#۶��b�q�����qQ��`�ם��~��#��r�H 7�{A���R��T�ɝ�mȊZ�lfZ����i�i��"������\E��#覰ʏ�چD�[��Wd)��c��p�D�����ӗ��ÛiT�n���\0�,��Q�����\���ixM謇�޻�P�j�=^1T�g��2x����̗�>���q���6r�\�z�0�\��g*��i�����E��M�e�����}��U����u��i��TTX��w�l�b�/�X�������Oc�bM2q������?�C�T�8�6��'��˴��
��b�� <�͗��K�u�{����-C�|��-�C�����h A��T���H-���-�f��'�_�
�=��&R��U��@�F��B>v�����{�ἴ��	��o�5�9D��Q�?����<�N��X�����@��?�z��HO��`Df�g�q�>���g����-ۃS��>-2D�6��3ꆛ�.���9����Jt%jqeM�ʁ�:���=��r:��`J{8s���`{�r%uX2�Y4"�巁�\<��Htބ����ŝ)�5*V�5A~{�߭�Dj�ʠ����-2�l)Pm@)�)������T�:��^�ϱMz� nkl�p�:/���������Na��Z�]�,Su[}f�g�!h�����B
�������@&}�͟���q{����a�<�A�ӝ�*��v��m�P	[��/�`�gcL��\O�i�Ղro���ڜ�P�v*�\�������͂/C�R��c��i���$e~Ǒt���O4�1���/����`?��F�5�8��@6��5���:�WМ�^8�¢��&Ņ|��SD��	��^8��Z#(#��j�R�x�$�b��[/��!����X%+)���?x��:�	��k~q�1��$��jzB�5�����%��͍��O�<)�sF��i�j���Ņ1+��:�1>$�A�%d{/B�ɚA�z��~��Da�h"@�U��9��� B�_�ޟ�����g�0N���8��f�jƷ!N�@�e䳣����`�d� ��h�-p��?4s�Z66g.�%2s���k9+���/;���zJ5�w^;A�7�&ǚ��c�`��ԉ�% ������ٜ���(J��:��j�K��s1��R�&�1��{�	��AN5���䏍&϶�ƈ��M��گ�_k��J�h>��'9<�s���O�P�5������p}����Ӊ��d]]9ʾbf�u�:L��j��d	�e`k��(�CFv�wIU�oWNd��`삅�W������c�p�	�9VϚ3�n�
y���1F�g�Yb@�A(�����	}����"K���f)*�B��:�f�_'�h䂣[M
���s+�A�p��c�s1����)����ޛg�C��� HO魁�)B��A5c˥�ԩ���HC`�s�R� `~�:�b��
�c+� α	`{iH��c�HUF���8�c�!j���ju[+���*��T�`�G� )�4��{WDͭ?z�2E΁NZ�8�&��<f��Lt
�&�	��[̧c�Etɬ1�`ύ�d��y���S2����&s��1s��1�0Ͼ96�� f�/��+��g�����~x�v��M_e͓����e��A׸!9R]@ ��_0�s�61�7C��1'<�slt���Q>5��S��)��4�Y�L�R��A����pT3�>���\�@B���-�8�f�|�3u-c$վ�4G5�u -��}S�A�������|��A�h5�;���Xx�J`��渐�� ǖ��c3\zz�5��	�&�=�tOwZ���UCݫ43����u����%�(����/A,�C��� �-�8Ǧ�ͦ�nt�E-!ȁ.uX�:��Mٺ&�7�8�%��s�{�9C��������ߖK��ñ5x �
g��<�Kd/��I�y�	d����)�O����Z�+�d�A����L��D�i�r�3�Y��QZ`��>	�4p8��fdV��V��������>\r�Jע��&1o�D`�9�N[�n-;��8�e��/��ͦ���[��[˴��G��u{'J�:�90.�g�?�	rk��M�-����L,�D� ��CW��ញi|'މ��[�هn�~L����R@ySc@���%��p͂/��Q�(�Gf��gw�H��Y�>|�oB�vMbvzM��?8�c�� n&����|#��t1�n{�Q>D�1c���ԡ���E�4�Tm�i��靵g��$���D]2:�3kWK?�o����C7����^��w@c�G�s��}Z⪧ұ��	��6�����(�-�����\#P'�f��G)I�(�rv;ܰ
d�A�ވ�I��1�ȝKT�p9���&��`_�)>��=�t�Bf���r��q6S�KK���=��8[�p3�IȪ ���?���"Y�P�̹����M�����|�|%y Oƚ3�E�R9
���7)-�e�2��������_U�� ��A�ٖ����}Z����?�!����*<�����p쉢�-9_'�8�ef�4��2pΧ���U)o1���vJ��>~�"Z��'��5-Q�|擭ҲTM������m)�A?IN����hJ/c|�/�̈́�h��vr&`�t�'�k.�..(O����)�g~���!����4��X��A?qT	 �V���ਲ���U%H��5_eɣ���ӻ���2<������6Ơ�*�[�O�aq1I����ꐔ��d���۝n	1[��;�е��sdP	I����K~���y}k��ޫ'��ѥRcrsp�yۼÛ���gw���plŷv�b��g� [g�0w��I�������[�����iR���u��0ʒ�,.���Wa��9��lX�p G%s��/��.W�)�5��s�UnB�w/�)A�{�m�C�mh4��{���T/PZ�_|b>S����-�02�h#�N��v<7��\`:٘��iԝݾ���0�;���3́�u_䒖\_��%��`�at�nF�k_��4��^xt+�i7D�9ا��E�����5��Aoѱ ����`�$�LW�ñex 7�-]~r;}_ӛ��/�]M/B�~�Yc�[_`i\����mqo�����F�̚������r+b婝L|Ɛ�h犍؞��7N���_���޾��a��}c�09���$���܌��:��qc{�IU����k�N�6�}ۖ���BZ�1��z���Yj]����޼d6_�V�s�H���ߑ�]|�̤�V-.�����z#����5ЫzK������/�8c� nF�aטч�4�����f�F���t��5��k9�����u(�5����[牣�U�w����m�4��]�O� �G��{25����&��?:�2���k,2-�C�r�?�w���iyG4Gjx 73�YČ�)s�(�߆}���<B)�fDS�f�2lt/-EE��<�*/2=�܉�+R�	�x�U��\�,9~�{SϪ���S䌾��
�.���gv����Q��&)����2*�A&s�Q��.N�Ѽ��jߒL�U��e� WeϨT)��ol\�R K]~r�(��1�9i�_��eNj�t�A�LHH�>k�XM�m֋~j���sиv��%Jk�e�N?�n��6�����8�&8N�"&!�-ie2{�,C&!y(Ti���U�IxDXXl��������>z%���߫^�ب�*T�Uvƍ"� �׷�"<���ub�&]���"�Z=���Ka��\ap��_���u`{݆�Ow�<E�tmZq��Q|W�%ev�.��f��{�(�˼��W)"�uPဓ�.�?L.`���E�V����<6v���[w�:�{t�v9U�ӊ8:畑eR����r���W�//=~(��?YIl�Yr@�r���f-븻o̡��-p,!�q��C���<5h���LĒy[�ѭ:�uv]�P��?�#Pd[pd+����s��@~�f#Nמ�<Z��A'G.aA�^�z��zL�on�q@���H'��K�����8M���N[�m4t��ol�Ӳw'�?\
�9_�3Mt��oڞ���3Mh���ĬA���q��'�������Ĺ�*AS�D�47O	X���b9GǋY�j{�p�c��UԫFK�#eu�g��cPZp������ӣ�1������~7&!��n�l[�U6����JK0�1�� ��A�������$�&:�jdD�)A�Wɛ��ǎky�����y�GG��|^���Ouݮ7�=7k�W���\��+�*IWQ��ڋQ��&m3yCr�����Q�Ts�p��Na�:?��A�m1�n7���9���^s�:�}��=�蝹$��Y�}l|I���?�e_*�%�����5�hd���_g��C6�!'9��	Wb��N	4��41�lD�V5=�����Ӄc5�""*\��;x����A7�G��Z�=�)_ؕ��-['m۝��L�~�i\�՜=z��sm��U�R�����=ҵ��L_�:P�W���O��szd��]��/-��?o��B ,��F�`J2�n�?�R�J,�I�@[����BR�q�7/�|����e��S<:8}�N��ށ��<[I��.E~�xp�6�z�F���L	[��N�r��8�ȇ����w�=R�8����8M�
�Y��9����+&ҩQKufaIAYx�3��̾�3�R Õ*ql�����w/1c1Mdp�+��+�Q�4ӊ�S��N�.S��[~<����R�|%tގ�>�3Nr��b41
y��>�k;��!q���JI�Տc"ö�o�`�<Q�`/b�w
�=I�#M䥍��.��Q�:��)!��"�?.=��ܿ�'C�C�Q���X���ְ�&��,���yO?��{o���5d�!Q��y��§�@�l�*��VJ,m}�u��B�V�y;ui��ϱ^�D����&Mjg�ߚ�<?��RJ�,K�"N#j�Q�_ph\��$�C\�d�!	�k�/<�s>᷃�V���ڠ�}p�|j���̈�ɐ��	��<�Yّ�g�4,�l^_O�9�y�R:~�
q8���]#�c���l�H��'$���K�B�j��I&�}i/�Dhd�\��P;�I�&uu�������l�C���a�9��L�l�-�<pA�;�����������O�p�wV�Ǌ���$�A��BqLL
.*�����99��^�zY�L2���%�N9V	��[�1���X,*E)v�7#�Z�R�d:��Y�ꔞ�]�,��7�z\��U�l:�����+~f�9�8B�V�х2���"�=D��#��[�����cX�d1$^A�4�D'$h��6�*�
྾��2i4д�v�/�l8�b�
��m����'�i($*��M�x��՛ݟ��uo�f#u����M�|̬R�b�H�du�@����Ϥ��ޑ~i�=���`3 ���B��h��C����SEWO����+A����RP�3z��z	b<�
	_$�;Sk
J�8�2��׷����
������8Y��%�pS+�	_vJ�X�Y%������忦�y�2�)�	��G7g�ӹ/\t��@{~�M��0:�Q���,��:�.<�E��Gї :�a�"բ+m�֣�m��C�z���:�9�q�S�=#uΚ��Dv$���nT�ɍ�E_=aA==���C$	��ҧ����pE��Q�DQ�]��E�P�a`���Tu&+�hּ���$������1U�ޛv�c���s���ޛgh��u��ƙ%�f�SZ�~|z �\���Ѩ��R�8Ȳ���F����a��ټ�<x����u{�0��R�3+��{r7]qw;E��B)�S�lC�`1W� .˪R5!�ȣv*����{ு��+k���1�B]��dSBY1����i�2��>`��ޑe�IA�/���S��5g��5��Q��D��_â���<$�֟�K�����������q���;�.��>�����"�-}�ccd�]J.���ŝ29{��x��2d����ņ�lؕ��*B?m[D�\3��_o_�>�����p�0u�sB���
��2Pˌ)�)��N��u/���[m_��ow��"�Նh���3��A�a��)�MŜg4�w�jzN��dÝ~�pQ��5nmd ��RO�ڪmFQ�K���|HC7͡}���>5[�����6��������s����r�^���z���1����4�y/Ӹ���%(����Sd�7^<`����Vɕ��=��Y��ʒǤ��`Aw��#:���:q�$%:6u��x�e�ƪȢ�K^>�W)x�l6�I�z��N� C���Nxo\�(����+l/��U+�`A��_v.�k"q�SP�,�S5UTWHNΆ�������HS2(T����1&�%5��#�m��\)��wN��s��-�l�4��yx��M˔rt5��a"��\���i�:�ۖ�ܿ��VKڻt +��e���/C�=dMa���vZ�uu�؈�[@e'w��ω#~�
w]?I+��Ĳ�� �LYjl
b,{�9-����q���㽹��;�0b�N�R�R��*���\����]9�NXX��i�!9I ��%$3�$[���k'/�?�������Z�-���H��U��}x�O������2��)V޸@9W����*Q��
N�iT��57�-ǵ,[��y��\a����$3�H�ݗ��T��?��YВ.cXGZ��^fRW��z ����,�rjAv���	Zx4���q�,�%����iP��X�!�@�F/=��}�s�/��"�l鍊��vpa��cS-d��8��rN.;��ZV�9�)�m5�y�����Ӥ~]
�����Ɉ�-J��M���� ^gD��\3��b�5<��(�����?p����ݪo{����_�����=]�i��#�v�Ͳsd�i��p�����A4�{�^iK�}�9��{+=y���l�;�����¢V���[�f�4~�BI&�D2�ԔY%��-ּE�E݉�?!�Q�VUq�8���Ӥ����ڏ�Y���ߜ���U�j��R�n����ݟ���;O��9!vL^����	~��ng���fؓ��7�wK��$���%��1-��P;��w�%������S����w�^�3)왢iHWq������s���� n.�:�5��h؅���&9>�u������4�p��-,Lw���"�QS��ŲE�W�����5)���ҏ���\!��� �O�<���TB��Ϗ>� ��[[�1ƣWn{{߂�N�+΢�Wz)�o(4��/^N:��X@�m���=�)I�݉d�<d$,ͤ���P��)[ArZ�:��o��q�H+����2����:XƝ����t�Vˤ���{�%�!�u4� �gw�D�=f������ڔ�k��FC�7KƱ��yJDƬd��R�
��y���n�)�}i8�I{)u���>b������sn�X�}��	���	ڷ$��d
��*U&g�e��@B]�ŭBIg��_���A����&�P���'+�E��(5d!'���a(3b/1��ݷ�8����[�:�mSm�V���	�]�C�Uo�\͜�f}>��Q8�����{I��@��$��`�[��ⱬ��#��Q���}��@F�&w��x�F''{ဤc1��9t�&����������:�v��Ԧ��}v��&�*�q,���At��Z���f�@��g�M�D��b]yj'���t>�m�%n8�M�i
�f���l�x���?	�(�s��.G���f��AW�~��Z��4�y����d���k���2�Q��~&�#;�'[Ɛ��) `\?��<��8��p��DR	|��D��C��v� n&��ݽ̂4��{?���4'n�<q`��L����l<{�Y�x�Nڂ��qAh˥�����%Q��f�@�<��}�z���f�9��t�[j�9��z��K���܌l�z��y��,=d�(�b���Q�I�"�["ZXLU��-���5�w�T�i��m�@A0��FG��-siѱ �{n!��{͔�<R�A���@��Js1�:�eZm\�Vk�=�
.���c�>���uF7��I�}7�Ҡ3�d&�z���)[.�?:�d�g��y��m����6�%М����3�}�N��Y�/�Xm�x��.̜�R¶���8�4�5�X�`�~�v��$|�k��`�#C��~^�8f�l3��e�Rer����������}��a�F���lb'��G_e͓�����P:��:���_�oZ��й>z�<���^�7"Bi�Gԉmיv_��!y�����y"c�Ӈ���_K	6�i� �.��o��ŁL<��Q�Y�9k<�~JpR;0纯���x�o�3�����c���/.�j�����i�g���5z~��߲��o_�:���I%(�/>Hk��M?��@#v���g
�]<�������X�T(�oW���f%�����~;��f�_��X9�õ�{�
5��JU�3�TV����a�X����u��<�s8�0��+h��-�C�64�N{�b�qD'7:<t�[;�V��M�D����*���@�\��F�q#k%ZX�?cG{ʤT��\IQ¿#`?���J��"��� ��HdQ'�Z���UnJ���l��P~[�s�-R��Eca��x��C˻�7j^�����Ђ�[h�Lǜc;<��b�6���1hH�x����r�q&���鰔Eץ�g	ryd���Յ��
\�V���g�9�8�c���c�����פ�:��(�-�<��_=F�7ζXp���~i�=��60��>���?�ñ<�s8>M�a�{�cR0+ޠhe�x�����f��aޣJ3&zc@��{�H
������ñ0��;��9`6�<�Z�C�w�u�Ѧ��ˁ[癞@jɗ1;��ޒ���'���S����-�ñ<<�s8i ������r:��M���{�(��~�5����cT�S��r��|�H&�聱�q�h���\���ICx ����󀏢��������)� �PB�*�0>�<;ؐ�����Ͽ�>�)AD��z�)�lߙ���;e7�df7����'����ٹs~��{�����s�+�p���f�Q*�Nh���pn��9�7/r���2.�y'�"%����^XMhU�[
V�X�7��a���י�@ *"��M�?���NB�VMp����>�-g��'U8�[	8�iEzCf�Vx姅�.� �+�iH����z������`�?�Oz���� �����w�: �� �w���j��+��}`��W�k\h�g�g�����q�P	B`A\`ZG7���}8��0����u9�l8��[B��cg"��]^���!CJ�gug%���kw�P�ݠ�=ܱp�*. ��J,�O�z���0���NF8����L�kq��ON��<�,�)k����w�z��ː/��°>�e <��	��s��؛|��ln��@ţ!�!._>=����=�կ.�n_�MaGں"܄9r�����09�3�Ӭ#�k�z6mm�6q�X�����fsaZ3�l��A��@ ��1m�oܛ9�s.�]�T���B$lL��-`l�\��{���L���7�#8o��'�p&T���^�$�.��������aG8��l���nᖀ��u��^�S7/�:z�+�@ 'D��G���{1I�7��Q���D/H|��1��z��;���q�jɎՂD�"Tp��tj���p�ݬ�����ɐ}��}��Z�E�A��(N�K�υ?��	�)�@ �8O�����7���~H��/��^���ωx�B�	�]=S��n_�b��������;�P���D-�_<io��,FN�s��A�8���ɽ�xX(;3����MEV3�PQ����'!!. 8��?�+�d�㤗un	?�]�� ��9��	�6�l��.�34\��p�j�cV#X]NTp�	oOD�D��1ūsW�N�@ |�J,��*4�k Z��pJ
r�d��H������0�DZ	�J�4��as1l,�׉�A �X?����*=HE"V�݁؎=tP�a��27���������������Q�;1�&tQ�B��]�J�K�?t7m(4Wi`I�U�X����圇�3F �@ ��Fr<YB()+A)�%�J�0�fCXz�*��@ e�F���H������p�/��U�e8�E$4�@ T_bjxi�⍡λ�tJ��S4����yI�������.g��A!�׎��d��O�n�!�7�C� �@ $��ËQ���<���s8r��棳E2�$,JBE�I�6�#y^1���i���q]�O[:��హ�{�r��4�ʻ���6�Ï��Z��8Lﮚ�&��9	���VR5Wib����W�%0>�.,�q�����@�>��t���
�gms!�8i5�����N��z��s�M2��T�a3�����嵳.8j4l;p#wڑowl/y��!��o��ݣ�&��W�2Z����K1������ߗv^懫֡ݺ�)C��5�塔���?^n�M;��@ B	ݵaPi�'
}�V�t���_K+'c��Uh�j�����B��K(	��k��Ϣۉ{>��ۃ��
���Z�����Fr��_*�v8w�\�y�����f��S�eǩ5�kH�߉��H�c2 Ò^8�@ �2紐�x�m�1��f�f���V.�Zʼ�p0>D�'�*}�����Y����g��۵��؎.�r��{;�����L���ɰ���!��2R3ΰ�	}����4�Cc!a���0<`.�@ p���{�3��QkQ���^�w	X���CQ��SJ$����1&���!{�������u'�SR{�#���b�,��H����3�f����]Wu�s�wT�'G'��㱣f���y�wW�l<W�K��I��m*��iq�#e.#[9?sz�OO�'S
2�npҌ�0o<�r�b�+y�c�;��J5��$���P����Mj��n�v�U*����4��Rc������J�J)�<�ց߲�� p�n�N�b��i)i݌'w#��c؃��LW�$^:�@ Tgj���\q�vm�����X��f�8Biہ ܠk�9�+ϧK�N70�J���sw�� N ՜R��e�Nz�P�Sࢱ�� �t�o��J�D�[Y+B�ys�� �H���1�ħ���@4�$�49\{����B��㘴��wdyq�W�������gbb�9�K v�悧c���@ ���-�Z�=jHy�]�KB�cw�lJJ�W!E��Y���"� .�S�v�v�w��66���1KRpBu�f]����M���#g]1����v֬q����˜�J�[d=�P� (��x�['DYr����cF'p�@�RF�5D�$l!������"��U�Rk�<T)z"T*�ɳgQ�^D��ӱ���P��E{�ȆR���J��	�Ȇ�@�P� ��ϚbZ" Q_�j�01!$�_�>��5XU_�p�ⱺ�p�A�@ �;9�3gs��&1�/Wt�1k�b��ե�Ĭ'��T-A j�d�9�L?I'~�C�T�@�(J����� >�9�KÔ2�i�N��\V�@ Top@�36ĩtéA�Y�2��|F�S�\+�󜎖)�#�&,\1?���+U��M�׾�Z�&Lk�v@���O������C��)�#=�g�չB�.P� dN��"0؂?I=�@�����Z�W��W��֍6e�w�=<9�8��L�Z��a�e�/X�����؄AM�����n��E.���!?9'��Z���<�6eP|[EH����������н�j��,҉6��;A��<E�l�oK�F��	�$���;�P���Xx�a�mƙ<	�N��*d3� Mȧ�&��JB�ک��aʠn�k��d���=��eb�A��T�N��iz���E�ϻ;ǭ���4p�c��r�C�}9��>t�"9aꊹ��yORr�k�U��JiT�5�
���V5���;�C�;0�Ԏ�}x+�v�&�M�d�vT'rI�O��G@-�=H���m�y��4���M�W��z��X�J�"����v��wl�WKI�R7�DiC�h����+��۪vc�SR�fȅ[�P�oܣI;���G&���
n��K'�b^��e'���Am����Xq$�mքuE�06����8�FgM�jJ_S3��̑ӆM���Q�)�aԓ�T}����I�����_<~����?nDM�9��T֞���/��6bA���ߺj�̾-7|�%����=f��"�g���b�:�}�363��,d�j���ƶ�B�Z�C�>�={����6���ka�xX�) �R�����+=F������(ʃ���w�k�nG���%�����;>�չ��%���[n�=޼���\�諾l<��3���׼�0��1�F�$���~���륞��������,��'(���9C_�����§����֖���ND�Yd3�0���֦Ah�,u�Gs���f8t]
?����c6@WM(�xHl���z�#>��5j�5���V���RR�E�I��d�0/֕�f4Vhj��{�@�İ���''M:p+7u�7[�N=S����L$��bن�"�d^�,���&�>79��ƿ?*��r�.�K!�EJe:e���&d��ϻ�������[���PI����G3h3���Ͱt�mU����ma��s1l:��h�z��C"�y��ض'��r�~�>��q�\e�,·�Wϖz�Ջ��N�V�|��2�����׋����A�f����׸G �b��|�$Ԡ��5�q���SPd5�Z��&Qu��ݦN�f�4���o{&��/u��-����f����-Xmֆ��ÔZ�A�!�6� 6U��mI13��߷�#=�CLb�X%��k�R��^p���V����gֶ��E��ɡ�Ž�~�JF#������*��htg��}��`;�����6�S���P�Xx��^�d���(!e���#ǹ��`��%?�:�~���5�h_�l~����r�n={��&��{��#�Mo~���&�=�Θț����WOOF�,���o��~��k$=Ȅ�a:w��׹s	w�6���fx�c`ٌ�����_�^�	�^V�m�#G[�����V��U����w[`l��ν�mp;iL;,�o�(�2���66��^?R I��B�>�c9�?�vL���7�����!P8�{m\��6ti�
�;���wCR|��)� �=��^:�����g��N�z�~�h�f<�lƔ ���Ҍ#�]L��ߢ���y�IЖ:z|�T=�Ϲȟ�D��'�9���
�0w�%�o\��?�.<Ѽ3������fP�l�{�l%[������]��=��^}��
'o^��L��	�ih�Q�o�1��ƥ��f���`���Bd]���!X	J��7�a�!��i��F�=�E�@؛���x6M�o�5��^���2J
O��P>��#��1W6�[v���.�<�	el6�`��6H�9�B���6$������p��	���T��A2ߍ�Ĭ>fH�e�`��3~��"H�Cs7���0���}�,t����m���"�!гi{���W����J�	��}!�}nIش�V������s�}�O �t������y~�����s�|�ag]���&l1@_mt��A)�<����i�2�V���� 6$�yH��;�p�f��hc������Y�<�/t�B����bg��aNx9]ǭ%�O�!�>x��ӫi<�yb۹���G/�Y��S�s{�3���q�x�M�o�i͸D,���=��{�W���ٌ��f`g���.x)]6y�� Vހ�
�D�h��)(��SВ������Z���BK��y9=��%�����0�yp�ϗų�6d`Y���L�W�@���h��si9Ey���I�Ǐ�\���aj�"�e�F\�������{���(ew~O�e�S���3��@��=FM�R`��壊ah��a3��[A'w���c3����V#�z�=���W����"��ߑUG�K��R�(IZ���z坞��%Q��~.ۧ��4r%�Kx�����_B��OrQ�*�����uJ�ê��z��_�y�c���Ȫ#�%$����b3|p��#-_3r�*�%�&�t-�ТVCn�Ê
&����n.��K�&���(�=N��h�Z�,�|t�8���v��'�x}�;Nݼ�?{��o�'	�G) !6�PQ����y��Բ���f�6�������!$pR<t��m�&e�_l�3׌c����VC��m�W��|6�汘��Zp���p��Zl��"qP8�D��S;L�Y=nf��ʞ�R���3)�_��8��o�wA����BQN�}�Nݺ���zm�\�yػ'Q)��v������}`B��P/�&o�~=�' �!�1�W��3QCe�)l��6CH����]R1�Y�׉��;|
9��Yv!�� �5N�0��_�s�����8n;�hι2��|� ��{���< �ں��y�����B.�7�x����9��w�d%8Z\ui�.�X�l����f�"� �[�pv p�(v^+�YD��] ����*e�W���1���q�<���K�_>L�t������@q2�n��`\���0�6�����¢?���l�B�j�/���\n.�4p��ӊ���йaK�����e|�#����,ٹ^yl8|8��"V�t7j%������}Fs��p㏜�����ln��r����`��q�z� �`\t�o��2wl��[7�n��Ϋqq�������!��sU�6�ۑwlKB5�� <��
�5�]�C�K��I�N�I�
͢��%�Q�{�����������^���o�F���Oفy���M�g��x'/�"�ݮ��.{@ˮ�Vþz2���znd�����Kf��B���]�o��Y�[����s��2�)�!���]����˛F�ػ.|�^�]��O����a7,�Z�
j����`�����P�����%6��mju�E��+�����5<�l�_��qt,?� ?���$L������29������\xi��S�����OmA;���U-:�����Oc�=�$$4a�)۫�X`���C�G�Zo��y�"8z��x�[
V^g,T��hdx^��c�B������S�A�'
^��Ŀ&p��8�����ӛn>s �ܲ
~=�g�����ȢBb��0}�&�Ax-n��F���H?����P%���b��}3��ٌs�n�/OO:��<xr���lٱYM�˾��x���r���'D�y��΅�vq�Y���W�g&e�[���'��]��-�vnH��՘iRK�}�0i��_n]�m�`�꯹�/O��6_���qn��ixHޅ*%�%�����_܆Q�\�u,�f{�F �l3��*�o��3�k[�K�,s�0��8��:�Mkױ�=���6�w����%K��@��	�y���E���&89f�H��n���G��'��]�5_�b�E[Ux�U�}����[u������l3~ɖ�L|���cGЮ�g�5OIj�!��x��mQ�Mb3*p����p�K�r%����G�'�,��Wyyc���U��ki��4�%��5�fw�K�@ ����,�ڌӷ%����������eʌ�-�9��I�S��k�f<j�)��QQ��W�q.d���9�o���g$��na-O�?���k�	-��q5��<A/w��^`!-j�A��xQ��w6�Yg�q)ó/���pj7��bP��Aƾ��X��،�B���mg��;ΠV�o�Umf$�x�����Tz�2��Ll�V�V�r��*;'�P���&��8�'��C6#%�?�]�Q!�eK��=�,���Aנ��i��|�S��C���i'LK�_�:"ytFґJI5#��U�-�Fu�mS����J�@p��6#����#*�fH3c{Gj؝��"��xh]��6��`�	�9��|=�]�Oߡ[�b�+]�����!���HN�&U�@(��mkӼ��6;���%^i��t���s^�d�����:4G6�$���b ��0Y�6������yExc�����M��jD��[VR�fo"U�@(A@�q�����'g6�����1t}�	��Qn�/V�����d��ؽW	@�,N�\Wt@%�7O׻�	8�:D �����i9pQP6c�%jX���!�6�>�Qn�����^���?���	�EHp���;b��4���SN�4�cv�(KvԊ��o36���Ou�8�D���i�hǧ�Nu�ͨD��I�4Hy��g\ �s�@��H^;�dH��Zյ]�S����m�m~�&�* ��E�ba_����j�|/'B���_��.ols1#���Ǐ4)�P�	�S� N `����'&)ols��zf7)�P�	�SN{�;/D��I�'�2N�Q�!�9v�Z�|4�2�F������6g� �D�d�1|�hAlFy!^Nb#����%��Y$ߢ?'#����f�EK!�)�K���%��"��N�"��$��0�0��S�� fJ±��4rEj�
�7lB�@��	��,��6c�����3����W��4.b3��r�����K\7�� �^,1Ej]E��>�0�lp6C��Y�V$.� �z��	xHEߏ�Dw����x9�
�_�g݆  �,�߳��^j�ɲB�E�l���#�g	*�Qa�^�jd3Ld)��/9����)6B`s��ox�<pBuF#s�.����06���Pω�pMXO�Ae�dY���P��p���Y��Y�`vV�<�J�<���T�1�K�;W�P��*��	�Rj��B�er�HA�w]��(pҐ�s�ꨵ�R�'ȕ�T^�ѩN�,p�a�@C-�@k��(���* ����+�ݽ��w��Q��V9�W%�����`٠���s�Jw�^I�ݠ��D�IDѨ�������?�FBq[=dȺjB�A�~=����U�pyu���𿉔��;m�?��]�S�UFT�:2%<���6�!�<<tw�:��&իڐm)��E�+�^y�wBX�J��
n��ו+�	]�!�vw�K����q�R��F'���*���r�!��DAi30\��GB�ҳ�DV�݁��j�C�y���o��鿥F;��@�� ��|���Pn9���!�s��*^���*=�WT�n��^�F����T����/^�9�q�o#.B�9��Y�
)�&��Up���U�
ԫ@ ���CwA-�X��޾�m��!!H�*6
���+���q�G�7����ȺBIy�s�^�@�BKn_����yVgb��x�_�������+g74�$�*\���59�xU��p%	A@���˶���d���̝zU�+~v�2	J/!=�j4�o��=l��Jü�&ⵔ���Ua�nRG��՚.����$N�㌻T��3nL�y�^e[�bO���Z�#�
:���Dtq�O��ܐ-B��6#Z��C�s�)(�������Z�F�	��rw��c���?�W���Κ��$\��RS뒤�j�=�3������T8 �l��^���p��!n<�ի˨^�v�%T <"�x�������Kd7N��n�˗@�h^6C�6cQV�>�S��L+��_��⍡΃+M�D�<Dz^w�'�i�=�a��Y�m��\,�
�ʢkH�:~I��7�A.�?�ni�ʣx	8&B�>�v�0F�]��-㌏��^�R�o1v[��q��r���V�%5¤�:�ԫ��3Ro��<�+!���
�sds9o�H$��D5�e�9��A�@����7��W����+�iu`>���>���r)^��P�/@ ی0=�o�o��?��y��������+Bo��$��R�n%���+xu���PD;N�.�*�xʷ#K^8�k]�s^%��G��j���NL��z��s�N�+�����J�ʓ;?��Ϣ����L_!D+16�L˚L�e��a����^��	���Ӊ�>!s~�&w�p�J*���R��S��?�Q��"
?�'-�c7����lqwN�Ԅ>�R9z�4-���z��wi6H��-���o^��� 6�&3�Q΁|��u���^�E�׫V�ћ����j���u�����ڦb?=F6ԣ=j4l�{+oʉ%����~��]���ЮW�w�?�[�YW��i�����AS�3+S3~*���6�]�aӆ$�W���S2�^�e*xDی�+\���б�3bNZ���p����G[+M��C9��n�h(Wy<^�8�fè���W�V����հ�C�ǫ�?�I�no.�����i*�@$]�A�!)c�������!�2q�Фx�~y(%�)4�㥣��z�$^���d _p�:��ٌ�9�Zt�>��^0f�vmm�~s�o���pn��'�h�m*�jAf���2?\��֍�:lL{����ԧ_���b�R\0d��<x���]��w���	=�X���<\��`����c޾�{`��5o%��%so���#a2������/I�vHy4q���Z��П �h���o��� ���N�S���슇���Mm2RW��L,���A-�u��5��c@H���`��o:l֣vsk�l���=�Yi�a�qjMvY�����g�k_]/��{ME�ȍ�l�$�f4����f4g��f\�78�W�J�W7v�1�).cA���j���m�$���)��d��y��x���lߢ7���r8�Ɇʷt�S�����N'{�b���t�Ż����]S��R�;5bꡱ�A��x0�&g^��{�]�Ѽ�y<�?7�U\rұ# �~�&�8���*����J-�f�:b2<��`���]��מ���v��i$҇��L��~�8�hL�z�ي{�G�J�H�8�<�_w}�f��稲�Ϯ�倾�^d��n�Xu����G6�+O�ѷ�#���[��9�x6��c��4q��[Ξ�R�qi��y\�X�]�-��kRה�^a�M2��&l�JB	z���2���[�sJ��;95an_}�,!��1kъ���+����u{t�×vՆ���x'��g��t^�[�q����x�!]�1+������Zҝ4�G�����xW��'sn�N�����ƹ;�ի@�f���y�wW��Y������&� �g�GL����z���ղ�M�d�ی.�� �ѱ�+]�q��~a՞G��YL_#��WѲ��ިK���6�I�#��͋�JmT�ٳN���~Ӕ�oד�J����9��\��_��Uc�]���x��W��+�( ���w9�3���yʄA'm U����.���^G��Ҏ�fT;"5U����E��E��a�R�De��dY�lW 8�������Ʒ�+�M��0~%�O�4Q�?���!�^���]/wE�'Xl3���o3z5�|���o<>*�/�7�׳���e��]�X�M�}fri�����ϰ�7��Ä��l����5�������}��  W��k>X�;Җ�-L����H��2�jK����%��9Rh[�_�;>?�Q�2���#NU�g����b{�j�$DY{�Jᴏ�IkJ�=ϯ�l����^�����Or_�F�ȃ�"1Ԓ��O��n�N��+��ݒ��̤Hк@%S=��<��ح{����zU�nՠ�p�>wȉ\	�.�v��m��ֶ����uS*�f,�l�HR+�!��wM
�|�j%Z���zu�nݹe��q�Ӿ�b
��t$D%mp�a���<�~�B�Y�v�x��
apڗ��Z8������c~<��-��p�K4���dM�S� ~�_�7���{��d��.���D���Y��)b�xU�#�an���@ .�
��t�Q��50�r�>����v���񰜷�c��H���b+�f�[�"fhKۦPU��LT)�K��P�S�dV�� n`�K�9�+o'�o�k`E�eX� C�<�[h$�]S��a�<n$�]�H��c;�dƵ��p�"�	,�	-�C1�.A&���"�)�wCa�Rba;l�CB}��<SK�-�,lbZ��v�+��R�חvU��f�����=���PL�0Ҍ>�M)I7- �����0 ��a�m����,�T�<%%��Ѽ�B�?�!�J.�@����O�ȷ��yf|�W	ou&!B\-F��ZNH3c{�chl����ֱ�q�K0�/w+�xƾBZ�=�Q����U{4�rQ`8l;�K���r	V��t�u�r��<�"�l���e>�lFO،EY-�na�C(��|�G�>S���� X�vI/	Q��ŲXs�9�+�5k�
.A�KX�8�ʽ��2��<Ěq��O��6%���

J��&N����N�o�g�>�w�m_lh������PC`�l�_;T�KJ��.h��U�ϑ0�X��v{,0�};J��7W���TV ��(�����:����T�6�)ꉏW�;��Z�}c���#��ZR+��m�'�y�/�uy<f�7A;AF��+F�r��~�V���ʜ�J����^}���WG�['DY2V��ӱb?�s�1J�Ԣ~��pi	���˝m3��k��ދT���'U6��֥!�޳�Mo�{���sM�'o2��� �I:B�#���w$66%r�~�Q��l��ԑ��l_ӱ�f�f,Ȋm_ە!����|�'�Q��NCp	%�^�q��*��Z_ֹ^	x�H�{�W	aR�p�K��P��iO�n�)����!)�54.�ލ���2�Z�hv��m�ӆ��SѲR�[vk�|ѷ	�FI	�F�z������$L"}
�R%N�X��J?��p	5��t�)�f��ͨߥ��c����Yْ��%6��i����ٌҴ ���A�/���p5B��A�5ČD> ��B��YO����;���I���ԗ)݆���p������&�ɿi�$�@`�������G��ʥ��[��Nr���޻pM�
�Y�d�}�%ԗA�'�Ss�(�I}�2.abBH�2y��eԗ*yG��5���v�g�C�>e������RU+p���b���:|?Rx���"����nps��'�I��\ɺ|�d�76��Y����om�Z5���r6��\n���W(:�5X�&�����o�h�T� ��-��ڛ�������t��G�
�&*�J���%!�2^�B#���/�?e5�4#ك,;��q�Ы1�%"��R�:L8ڞA�|f̕F��E��<���)2Ҭ�A�K.�XM�����w�"����pF���l�J�������������j^
8`D���=�3�O9�.�2E���3˳�،�1���2ah�=�1�l�T��$�6B�F������~�����N�L\���}�lR�L�ר[�Z�F����2�j�1q!@����W����ҿc��w���Si���2ltYY�<�8-qP�Z7���~w����E&@M���܁DZ�apLQ�Y��p=�/��I��
��JL��>7+�"�O�:xXk�v	mU��A���֦W��æ���N�/���b�1vE�������lp+��8�~d¤���;�X�>5���*m_�6*�[E��/[�`��9z������mU��:7���#����`�&�z����iC��Si�b�<���Y}ϸ4p��D|�x�9���G8��E�9�
r�D�A���:8�S._O�<����4O�*���
[�<���]���\�5�e2q�ܿ��j׋mƘ�u��"b3|���B\ҚQJ$��:u;e�8�Fy��9���!��Ųe=��v���)�nO����-��gʐq�i��DPr�ŷ�(�#�Ѝ�i	�~��9ۛ�����N�&daiCk�~>����0w�
f���8Й�A�%u	4B()�M�Y��8=mn�<oޓ��8��Z7;��ry�q�3lɧ%NK����S�fīu)jd� Ȩj����A6cV5�3~�T������6<�~N�T&}D�S6%�_S3?�̧�ޏW���e��#S(��K'|n��~x����Ѩ��GE;��S�6���:���t�y��m�y"�싴���Ճ������\9=F��UZy��&8`���ě6�!L�
��,��j�n�\�������6ln��G�y�fu[��f%��ż\W"On�P{N0��GO]Xj���z��1��W?G�Q��W�Qꩍ*ω����v������6�?�f,���8e��ѻj�<&6��^!�M=��:;O^�ιq�9��p�_�/UMk(WG��{GJ�TbX���&?���[�v}���溩�{��P���&���"��0�}lv:�O]`u:"�
�($���i�e��|�w� �zg�j�0��ob*W&�'�0q���F
5�Wj�^5Hy���r�וbq(�W�� 쁖Fc��Fc��]��RF��e������$����V5��x�
ڌ,d3&�����]�U�Z�q�a{c��h����}�1eT���X`EJ�$$����%:��+ܡn�շA������`�_�;]7�� ~��c��P�
G���}4�3_�^�"?o��K�V�Џ^�ZV���cr����^�%�0�gTpU-���+U�z�g3�����D6� ���/s/���,�D*F�e����-5J�pԷ��p�x���x_����S?���CL�Rg�eE�8�ڛ����_@ Tu��f�����imb ڌKv+'�/ըϥf�Z�q��or��M:0[����Z�n��0�����q���0s������@������6XmƬ?Ԑ�W�ڌ363,ʹ /DՅ�R�fC�%A)���Ey��(�>t��ʶ�R��b�����O��q����s��mN Te����허��%�� �<��޺�D��Z
*79ΓpSq>7�L��"�>�|}IHp���~�rkU	��)�ߍ,�>���ہ8���4]P����[��� ��#��&��J��5�����X�A=�Jv��	v����4䠖��	��-\�;X��bO,������P#��^��i4��!�d��@�T���oI�>��Iï7 ��&�(��m��
��JqzOP���f�rݯ��2��y�-��/�����XsR�.ʸ9.쬢�*���ܼ��g*��P�P�)�3�`7(�f��s6U��;�8������T�=��J�M��p��t���G,�W���49D��~%,ܢ
����~��xw���&6��A���ms��>ߥ����`����~=�ޫR.����r(����@Jl�g�f�Ï6c�5)7LNlF�@<@ȷ��ӝ*nk������J�:4��K�|�A��c�Q��ʟ�!����<���8;�F6���6c��!�S��\� 'r)�¦�V�Z��#�ihW���N�E��8����3�B?�/A���Qp�:;/K�9+�P�8y�~�ѭ��g3.H�d��qٌ�f<	�XDnX av���x{����
)��0:�`����/��d�@#�R�*^���b���ej%�T&��C�w�/��ǹ����4����ݭ�~�f���(&6#Hx��}�=B.E�A~���d(�E�<m7o10̧���,H�;kpf�8�1xh�D�F3�����V�����g��ͅ��_����{�����S�7�*4=B$T��^��q����2��O3�W�{��C��Hd�7U��+�V��K9 6#�a\��_`JĲ� �.yI)�7«��A�,#%8��>SѮNs����o?t2���&���}j�ȆUF'MH71g�w���^S��N6q_jF�C'��]���v}���JmFgMH�`�^|�w\��ö,^���	�z3`�*�ת��I���gvT�t�����+���E�(V$:���]!1���uӘ�� �ƺ`�!~ւ�iޜ�~;�#��	szhC�����X�N�l���v����9�Gswt+��0��>lJ�%s�ɋ��fg�_3ӛ�7~���v]�]�K��B\�K p0���tu��5�P��k�l߷8�vHD��F�9'8c�@X�ߖ��O��{Y=?s�s�`� }�w�����<m1�/�V��emj�T��!�A!Q��z���?�V��eMj�dt���At��:y���^�k(�˹D�� ������s��Fa;W���ꖓyqB���\t2+5kBE߿.uͻ���tц�� `�������ߩ���/X=1*yx����f�5˜��튾�7|�3F��	��%TsX�ڵ��m�.�8hF��:0}ٍ���v�@�}#'g{��k�r��Y��XT
�,Pb ^ ^B�A�d�]Cw�,C�2�����E�q*�Q��r�NI��E0ٯ�P����:������[�ǩt�����q%�����/�}�'����C�p���H�`�c��>��a݉�\ϺQ���g�oݼ��+�%�XX�x *��sF��{?]��g��|ә��$\�ᶗf��B�ݭ��E�9��т���������|7�r����eV�# ��xA���_m>��3�}��x�w�^���l��?��@�,�ט���w����Ls�&�?]h7�@&��G�ݱT��
�o �p�B����2�ߢ�\`��6����N���K ����p<��p�s��m�(�$�؉�d�@*���+�?C�8E��U�L!ǿ]@��u�$TY�p������)����!���9�;pj1$5ZV�P����H��@gu�5,],�~N�p���|N����:�KSb��k�X@��Y���n�?�:ò��O6��s~�0��)���E�)cX���XУ���wp�ά����c��.�3�%=��b]V�E<����������x�d鐙mx���7�C �;    IEND�B`�PK
     Y�#\��ZO%u  %u  /   images/c73ef27d-6394-4828-a75f-205a980bbd83.png�PNG

   IHDR   d   �   ��z   	pHYs  \F  \F�CA  t�IDATx��}`TU��ymj&��@����T�����go�kYw����X��P�.
(��tQzM�@z���y�?羙d2�	!���d�w߽��S���Ep g �џ��g?~��g~R��n�)��cg��߃���7��� �����s1~�N�8v���
��B��]]H�&� ?7�gd��	�g�m���e��o ���V�u���Y�����u`QU��Ѹ��tAC��#]F������Yg̀��\��b�������+�,�
C�~t��2 �L]���	�(�>u%t��4�&�Aw�.'���� �{��.{�3���&�.�7�x���8��K?�e{6AW���r3�y�bd�$�[=� i�p�ZeR����頨���M �<5TZ�}�_-� q��bx���UƤ�������=N��G/GUl]V�	�Lo�W��������2������������)�=��|A��m��H����f��E�"O9XU��g��2Z׎��x��*NR զ2��	��J ��������)���@�>��UaCԪ������ȈU!JyȮ�������-Fռ`w�*��xN�Ds4;C�N�Îx]��H�9��R�IN�j�2�Ӣ~����\��7Z���&Јp�F.�=����9U�z��.�}����`bV��󈃼Z>�f���[�ގT#!\�E����h�n�y͢�g��O��0M����>�w:�UE�&��b�3	;6��>��F��5��MU��x۸��]���u���uϣM�1�X4���`��!D��1�C��GI��Yv�p���"�Ka���	E�5��`�%���B�a�oQM�|b����n�����NEy�A�͍�Q����+r�/�(ӆ� �.;l/�&_
�e���z�L�A��!9�7SH���~�h7|&hp�cAV�����A�%�g����#<����q���e
id/|�8��v,�-C�x�q= qXV-{o�+�hQ���O߭*�j���E#�^K�$���Y�OSם����5%�9T�f����@�8��H؞�_,���퐙�L���T���),�n0�pZ�I{�(j=��8��F���J+��m��\�T��'�G�p\��2���^���1f�A��MP|�E�p�.�$�ESF��p���F\.v!����Բ�ʙ(�&�=*h�ZY��*H�"�5(�dhi�*5�<��Q�E�{Ks�7R���Lf���;m�pK��:��9<%eԲ�V?MV~2�Z&��;Nr�{�����,��F���H}��e.wo�0cP�rH��X;��O����\e��$.ơ��R��F�'��W�d��y��G߃}/����N2Q���#*pU����:���(��xyX�d���|h�N�=Y�?��x�9�D�>�;�#���w���Á�:d�h�
�섾
�vr���i_P7��+p���l#t;@��^^��>��P�����&(�l�?�j�F�n���'����������1Q���A^ؒgh[nE�,��l	T�<;e��ƚk,�8%�J�}� �P�r=,�	�����8I�����/�;��2|R�m�� �,}���Hz֫p�Gq�|��9U"<p���Wk��j���D�Z��D�g,��O��'+�Wi�r�8�V&XT��.���n{y���&6h(7m1�i��a�rK݈/@��
R�Ps��8Qj@|���,�%A��e;W\.{�ºJY��&K+`��'���ہ&��x���R��Q���|(t���hԻ�&b\:ul�5 rky��4�����?(<��:����Q:���ԖֆO`�&�**�s�y��~����5�s�9Y��*Z�I�4~7��+9p _/σ~&++�1��`'�����o�Hb��x��":����s.02�_������ʻ�o�K�Oq�Vn ��?�~߲�?ěU�6j=%AK
���pV!�h4�?�k�ndH4�\u�Eh���a�
���7�o�AF��S&g���5��Oe4.?�����4�@���X��a���: ,�
7�+�r��_�q6�PZ��] &*�2�K)��t`�ϓ����Wm�Kj�<֬}�>O���L��Xڲ��>�/�+����5]�ho)u�6�����j��ۻwlٲ����x�С�`2� 1!����T`{�۹k/�ޝ͞ML���Hd�$Abb|ˇ�O[�o�G���Q��	I���ѩ�2�^!�/���%��;��D�������[�97���Y�� ���ĩ�f@9�z��w͜P�54�����ufiN��0r���(V�3��rQ�A���/�\k�mI�jeV8�-����$L�v�u�M�ӭ���7o�w�j�/l!,�*�~�&X���2y"�{�����ا=e"�|� g�0Im��(/ʟ_m��e������j�0?��$��ųP72\,��lauD�t��Ĳ��������ћ�PJ�Rl��
�:����s���퓍�6��]�c_ne&e�WK�����r*�.��B���� �"���"�]�� �H�ѳ$�@��qq1�Ђ�A��y�'+L���u��&�Ss/i����_����챍��N�9�i��$��g3E�fo/�}&+)�U�����	OD�;�0��{�9t$c筒6�Ɂ�Q7�W��޶��sa;���p���B||,,^���U���#^'(�>��y_U�5�{0�8H�]p�YL���u��냔�$��9��i�Na�4�Fx������-���74���0ԕ�hDM��#G����"."Ƴ��I#��cY\�(��F��'ld�ʚ�mv�×�%hIQ�J�{"JMuߢ(ȫ���: 1F� �T#؇b�/��`�c�D#�~��g¤I'��%�aٲU�F�q<#@C��I��(��7�,+���g�uC~uUpHj�d2�y���%%%�������P����saP9�8���c#�xj���''�1j-+rH/H8#.K�	�1 r�ޜQMŧ4u�	�#�O6���	?�xa�t[������:�ݳ��v�0��^Ye����p�HLCVO�)8[92w�����3��E!�����h��+���,� +� <��S !��Tׂ�|�ؒ�55���?f3�WUU��mx�^���s���/Eq�f�ԇf���e���\�^���<����G�T��q5�/v�ڌ��F���
؉~Z�%��ۋ�Cqu)��ԋÚ:�wO���j慛�so0�у_���>JQ�����dɰ��D7x5������ӇvP,k�CU2�X����^��7r
�9aG~����UX�����)�B3ƈ"Q��}*^7K����H��	K�zEi%��� aLL�②8�������Ę8֦�K-R�h��������W3�2J��*6Q�Zŉ!��[�9v��EcO���
�l�����/a4ȩ*/ >�X���F���]'8�6~�ܵ��V� �}s���77�ё�C�gC���EV����u�B��SQ��d ��s�}��ٚ���`�N+lcy�/�� �9l d�w7-�W�$�&("}K�N(K#���#[�W��� y�� +������>V(�'����4tAw�\N;�l�M�*���$�)8�x+��u�k�钒\��7�H%�Uh�������M��i���7�wٿ�āi�}�Q�(H�'Ͻ� g����؍�/��G��\W5Ĉ��]�>3v���\�;wW���,vg�GYZ�L�L���AI�VX�lS���-'X�fZ"9%.}	<�7��@Q���O���x�pRT�}%^�/܎�(�.�
��@��hQ|j}�#� Q��ٟ��(����4R<���n�_[Fo�w�-!B��oU�&x��0>�$x*�E|O� �m�h���@� ^�?�
ؽ.p�������� B�koY�N磘O��,��-%נ���d-	�Mc��g��_\I}��h���9.�F�A��Q��������	�Laz�Wu��t����W7'�͇v�뽈�Z�#��p�C�셗����/Ji�3[Ųh����*�;��JD�#���!�,!�S��7>� �dT�"[e�����=2���%O8���������%n�wa'��6cYv��	=�u�=๥����M�W�z�^�Y�a���vp.YkH���<#~]Q<�j���1�e�D��C�Ȝ��0��>��$���	񿋽�>��-��Z��Љ��^AC	at���D��jG��'D�)CN�_s��ӭ@ZR*\��xI}|�s-L�3F� UȮ��ZN��c�?�?��'f���m��&�)�	���O#&C5���5p�Љ�71��`��_Z��D���J{pKj��9^h0��yY�['�U�%���@T���P�7@�-��b᷼=���������VD\<s(�ظ�â�L�Q���ٛaL� X��+��Sc���[�2����>��9�̡��w5�I�bX��&���Ȫ�⅒�ȥ�m�5L���U�g�%�=[��5NR�����Lpz���v��dQؑ+{=:K��/=����W�A��t�@�(����NF��&����^t���]=��O�Ǒ��uL��;��S��9�o]�O��¤�]T�@]�z.���э����|�����Ig�g�(Qai���pf^3�lX��j���a�8S�¡����1���ܲ`��r��-	U�z�ی�O�
Ŏ�B�0��VEc�6�b�_^ ����0�G������5@z|
Ԡ���P &͔ uU5 ���(q�걹N����()GS�5m���o2��u��ī����$�J�G_� I2lB�b�]�����?��k J�ֻU%�􏰓���E`F���B�?}
"�����]��5�6Å'P+�<|&,y�t��l���kΆ�]� �<(D��d�R�����3�WXS���Y8GV|��֕`����b��	m5Y�~3���ع�B��;.�g����������/F��ȯ�ˣlx���GI?��A5���o��;E���On8����
U�̹V�b&�C+��#,��r���u���$�9߶X�ًΨF�Dr���.GS[$�w�j�����+�B�|�:;F�5�[�B\��D�j^We�m.G�-Gq�"�ǋ�È���;�e�s�/|㩯��+3{Hƻ��6m��A��)6��v�ה��&�q���e����fe3����P!�#pwd߃~�������0������=�<^�1!L gH��*d��7��*���\h��iM�B��x���ŏ��&�ee�t�h��ޘ}c���K����׀umj&���\��sKA������8A��kiH�٭
�� LY����(,̈́�m(oV�Lj΀��
���<�卧o,�	ߟ��A���wyF��͊�^n�U����J  �Q��WmcK��84A��&�4���qpЙ�*��(ꐻF�?�]�:�����͂O�ۡ���}Q�� �C�;���Cx��:�Ն���W8���0�:�����U�x�XJg:`;*���+���bY��N�Ù���z��Y{C2V�����H1����S ���>c�ɩ�¯�?G�����c	�?n�e���a[�H�8���aC'sd���+�+ᰠ�ܹ�,�;�6���2e#�h�յ������|��$��dcz竪-P&Ww�@^>�$1IpH4����r�XZf��&洆�x���!od�l��Љ��  ]�ߒ\0��.��~/��T�"37sD���β�8=���PXU�Z��$�~��$�㰚��#���B�W��o��$����q�	{� �u鱬4�E�hjX��YC)�GN�cg��.�Ґ�h�Dҋ2�x�R�dR���I։Ibg]c����m��yFaD�*ܑp���0���Vْ��%-M�D��]�����|Z��͵	����S�A3.��l�۩;�70Ϝ�g��ACSI(��.��흎��Ѓ�f6���7x~V��WӲp��&��5�7;Q2�Gۃ)y$����/�'5�g��!ˤ����j���6�U㑽��T?� H��0��fxk�ܠ�y_�Ԕvj"��w$i^���N�������~[%�N��)!#�E�}�hG����A�m:�ӻ���g��;4_�F�R5�,9V�iYk�@&]�ꟳ�L���~�Ǚ��S���4�֒�V��H��
}������!��G83�;�RV=�?���B�0_��]����_Ј������?�=s�]��(��w;f��W��V&6G�r�M�$�UpgT�gL�`�㈞��=��d��@Z�6���C�k�
����)m�J��А(�3�o��� �L�h��s��P��ZaΊ�na�ݚ�/y��
���bS^�>��z�я�_�}�n�ㆵ����T]���f�sT�J�7u>�r[�Dr�����Z�O�s�u@���U�@�#'��<nT|��B"�E�[�(����4(�T�M8�4Gs�&�����T 9���ɓG�o�C�����T�x"�r����d�0"�� �(=���/���jG���H�Qc�&��&T#R6��>P����S�(-J��2.}��s�-�k��O`��*ˡ��H̿d�R��0�� ��Ʌ�b����=۾��і2D�����ˡim?����A�/����	Q��	�!5�����
ny��R�9��Kڎe�eETD���b�Ĩ�Ѐ�tX�k�|�6�`�Љl���,�`���@�x<PWWǢ��IiM͎��P���ˁ���,���|O�ǲб�v�vIDZ�e�(l�_N�������n�!E`�EA|b���B~~>���3B)j�DٺvRwr,�Ӈ�	IL��sF��xPZQFǈAȎqqqlO%5)j�QB��b�M)��^GP��}G¾�|�s�%L����[=������^�q���f�ACC�۷\��_��Z�h `Y���l��)�f)>j;�aѨN��R}�1��FCMc-��Z��� 11�k��n�{�	O��.h�H"'^&�Jj��Cv�_��}Mc5��-�^<e�x�~�zF�Ʀ��ŉ,K��O[�F���F'�4�X#/�I��!I4����9�w�U������ɢaܕ�=o�LٵՑ9�O	q���n)�P��~��!�_�p�<U�@B\��S���^M�����9-�6YS�ݠ�B����e��ɰ����4m�����'�bɒ�Q-ZMӣ��`���N�*�sGN�l4w�!$��(:�3<(��{��{�B�-�Ab
qG��oĈ�=�����_O�N؂9;��6#�A�}�؀�"y'�����߯�\���x�".�K�H�f����qj��'�� �le{�@O���CAr�8U��ڤ�B_����p)tBn��J h�3}��͔�]m�٣������'��ԩ��"_E<��:���O������J������Q�m	����l�*�|�����+������4�r��B��a��f"B(���v�"�RD����w
�0µ��c8+E�x�)��u���H�>�cb�(Mn��ͼp�9=��;|��q�t�2���`���W�}�d��B�c�����p?KĶ�����!��B'��B�����,�$�u���u�$
���\oL<�>�$�g��;R�LG\nE���0O�	����ʊŃ�rr�ˮ���oi&Ų6��Z��@��/��QS!E\ZWcz�w�-�@�'��J�Ey�ZgVF�6(�\4x"��T���Y@H'	����v����0�`�
�,��p�-n@�h����A�腑x�r��T�:�*�DД66m�#���%#>�Y�-��:���� �b�:{f 9yQѶv�����:E�!zǧ���΀�K"}|�b�'��h�)�΄U{!���S���N���"��o�N�X,K����O=��j[�~x茫Y�{AM9#��،������67�bZ��/��,T���.{��nh9�K���`�|h{�~Cgǲ~=�v!k��g�,��f�= ::�����m�"ill�>}��d���V��9�u�S�B�g(K�����
8f�L���$F���
HNN�����J�$o=!6ο���X��֜��9%�r�����X(��{*đ�p�ẓ΁��.`y���C������@Yi)ؿ����l��T����Am]-8�ׯ�Vg^I���ʮ?i�=|xQc�C�L4���}[�����հ�DP�+�<��G���E��{o�qD��P�h`^���\H��e+�2�eՕPQS�2��a#O�SѨ��f�߷�C���ч�im�$Ilk����|�D�2���
�u��Db�Ǳ�����O�0+�G�,��%n9.%���m�U��D�0�d�U���W��F"
"�׼���̫�b�.�Gb�3=B[�f�� $���ﵕD�!��"Ze;ڂ؇<�p�ݲJ�OZh��6�����G(��@��_��mqp}R:ED>��6��.�8~B�m���{9�=	��ٻ.^4,�/��u6�9�l�IC}P�uyfD'޸	�F@$��ߖ�v@1#�9�lq�}T���~c���N����_�ϡ�B��`|g���Wj𣏕�3b�V�{=�����p|8��q��3 ���D��.��F4Lk�t\vO�N�����`�5�Q,k�Mo4�ˢY������i-�����6l���]��69�;�?4��a�E�e��Eb<����ŷ�T��~A�6҆P���y>�e!�������}�M{n9�M|���+
�pmƲPd�6x[�*��f�![�Y��k��H@�eU"��-�}���߾�&%��8<I4��|$y����;b��,Fq5���H��&����[�ր1]�2�����Z[&��bC�W��0U��3���)��~k�������o� i�j��u�X��g7҆����Q9���F	���7-�($��A��:\��;[�1���mL
]������Sz���Ƌ�X=�
�ޫ�-~+{�{+�����o��Ų8���`�\^�8~w�"��&�{�^��+����u�0����xp�L΄��BX������9�Пy(�7��׼P���Sr�Ԉ?�ޞ��n����9&��|!ڢP騃�7.B�P�A��F��Fv�H�/�`S�^����iB��z�p�X�j�" ����������W���?Z��"���;	r�M�&�i����_AN]9�6ԃ���<������~1�j;��� ���M� G��5�U8��$(��V�,,�;��|����u�R}y��_g�hʫND�Z���IZ��v� ��2%L���Tx��#�*�]��6��ye�1���`�R�� ��֚�Յ]���HF��G�pV���Ų� =�� �^���I� ����ŷ���o���vY����-R�Gy��pN��}�,�,�$F!��%q)�D�p�J4��L�"� kZ~�L#����y�� ��rǐ�1Á+= �d�;ls� �zm�^�"W,ܻ�Y�To8����w�P68�7'gP��b���9��	�MѴz��~.���R�,�_Ų��=��Fs�D[�o����ؤ+v8:՟pv��<�N˹�*�D��oC��F�D��E|v�-��5��p��z��Ѽ�ҋ�?����d���XΖ-��O!�n��lk�)���0�s`+��4V���-�mnk��-�`W���|ٛ�;��뮁�	���
�"ܵܵ�]h�8:�W��̋��ǿ���
�Љ�����l�R��`y��b��
��� 1P����l��j����3F�E{/(A��uD�{
u߄������q��t�4�>F��CRF/�*>�p(�up�XE;z��N���7A�ϝ�*�&4�	F�;������Ҵ�ѝ���d�Td�>M[�VQ�0��K�*�W�L:NF0Ml���t2%�J���$.�8��߿��</4p��I�:�w��d\�VQ�Jl7+�`>��Eb���,�%�h�UNd�0VV_���8ShŐ��^���BL&��:*��Z�2p+^�y��F"X،`�XJ��S<��}��	��9��?eyde����5�mT<��W�_�<νe����"��Gd]Iص>�j@�	�1F&�$r�S��D���-�v���Q?���&��mMj����W��p[7�o�o�+�8� "�@[׺��z��ɮ��X4�J�Ϸ�tl9����Q��iBY�<���e4�K�Cm�M���/��QD�cY��N��d���3*���/k���� ���t	$oؽ欢C�&�?��6}L����vNu*^�6�B��1�?�ԧ��6���f�$�efJf+�%��|�����(�J��\�"�#X�&g��Ğ�͇��JT%1���&���B��i�]���`���'ב���T;�G#���p6�d���)t��iY胜��^F0�*�oT�Qwi��{m�(}�*/�OK3�rn��x��� q.8"��/Ӥ��;.�q�@8���CU�s��^��	(�������ɉtO��-�d�H,@GHQ�oCbY���r�2�wŲ����{�#!�<!}0ԡ�d��M�5�נـվ���cp���َu9>�ox�\ЯW#�,�E\�I�D��i!��Q���);6���D�W�L�#0�ԁ��A4� �8��G�W��a����M+���J�4ZF.�Q-L��oE/h�ĉ�U"�|ʸ��&�O^U]�����ސZ�mϳ-��.��8s������v�o\��mG��P�qx�~���`�5�d�E8�i0ף���v�����۲]n�gD��F�>ݪ�����;��@����U������?�Y����(g��u��TXM��ii:q\�Y�lœ���:���n��+��A'T��Z�1��x�Ш�R��Y:"�×L*Ń��-~�s����DlP:���";�ڣL�vI�|>����h�FA��������4H���޲\֧a=�B%�\]C����`�mE�Y�����p����j�%`����%��h\4|�4rj�����m�3��I�7�h�׷,�����)}&��FA��^۳�E!q>$��a~�FXS�3l�Lr(��&0E�����#ǐv�jjg�dlԞ$A]�D�w;@���o�%��^1lU"�U�*\�>���5T2f��)�}�^x��F5�Bo�]I#L�L����0�d�} ��ΐg�W����8�I�$ ���P��r���0%I��-��jȱ���,�d�ܯ@t(P��r��?9,n�?�6ǲ:Q�"k�,���Af/������n���
<v��4��P[W�*��]��z���CqY1|�y/T��ːxVX�DL`Kq��SB\���o$�L�h��*�24���I����� (�uL�������ȿFd�b��gj_�����5b�+ͅ�ÇA�l�oă���N�L�P��� 44'1�ɨ��d�\��y2d��9{�{�U����'�砃%Ý��z�e������2ɢ��H�#U��Aڂ��F���\�c�����:�\>�e��(�z��D˿��T�tT֖�zp��K��ѱ}�B,%��� T���#��S�A��^�["��K�>6XP��T�i� s 8rn/�1�D�ejrF��Q�����k����Q!�mC���`oS૭��%V�dVآ����r�l�Rfe�x��d�a�t�"��m�� ő�/�Ͽ�ű޵f��N�
��pvyK�xc�^���~�z�ES�l�6Os����09*D��Л��f��ǫ1������2�@�\%k����h��FEW��8KTF�g���8Tz�z�Χ�47c��u��u��m�.���^?���jE:���҄.�Z�Z�=a��g����} Jv�4��T���oC|˲E]%�
�����;���@�(�jP���h��NE�ᦤ�E�Ŧ�|ɝ�2b�1pń����
�����o�N-M�Yf�@��v�˵c��;?��y��7��ϻ-������(V�e�/�Р��i�}]܍�)��h�Il�݀jj�`K��+7��9#'y=��I�d�i	������{J���؁���?����-oO�l�3��k�w�vIȠ�}X=/+�g��~rubO�-;�O�L�^��l�����5nE�t3�+1N)�8�����cȊ���GN��NV��L�!���!����E��-b��)�A�%��%+00%n�?
j�&��j���(?۶��`��E,v������g�pF������'�� +�*cFXc�4�q"ύ��墢�?�EíbPZ6��~c,�%��U�w����ө���IQ������i1�l�ςU$��*@�46!�kK�b�i�n�n�q�Qj��c�d�G�;Я�Zp�G��pF��6���!.%li�記�E��D~i�[Q�� O9�	R[��'�ayYa��#���ϟ		�բ}��Jr8�߻� �u�>샲�0�i�"��.�8!?���a�}�&�~��Z&�;Xaq�Kc)m���P��C���p�jO�_�����R8|P��63i���Kf1��o���`_AM)̡�` ͩ��I2�h�5"�,HkrA��x�	�©8���"Hp���⣫�寂񛽎�nZ_g���=��<�Ӵ&;<|�a�IC��q��/�v�o������P�Cau��~��j��l���`0EA����A�5TAr����v���_���;"<�R-��
�!��{O����uEH�A����

+��Ơ�9{ЉpEt,���@:κ{�,���!'jv��|��| @^��ۏ���t����ͧ��8�>��=X�Gμ��,���8�v���&hh��XnT�k�x�,N�m	B��n`�%�œ((+b�\�5��GkG�w,V�3��U0�Ik����V���qP^[���!:�WC�=�D��[���ڲ��E�#�,�Dg�N���D$��z�J��{�����M��H���A�L�`���K=�T��PUҍ����Ue@�~�m��\�(��{~�\]�m�2�xj?�����
��\@ШΕ�+�����vAu��s؏t�'FŲX�a�%>Z1�ya�7�QZ8;i��}���3_/χB�3<��%�Q7{�!��%��%�7��  ���(տq���z��;��hFߑқ��s�y��	�����,�����E�	���	�A���Z�w�@SԺ���㭱�͊O��j)?,} ���X�E��[��xg�B���Kv�"�`����?A$���CbL�������;J�[�f�y3b����쓑8K�0�f.��Q�yh����;h�T��(A�k |��X3�d]�YUL�N�sk����i��j����N���j�V�09~ϩ����c�g:2�D}iAH��$�����f"�f4�6�J�W$"�!������mu�#N���s]�ϳV �l��bYNEy��� "g@�棸Jt��=�AE��ԘDw<"�7��!��|���{A1�I4���uG���m �EY#n��#��((P�F��./�)t���EVS՟��mHK�e���������E����#��/���ۑ}�"��8rN\�t?Fb�5���kБ�Ü�������f�e�PI���Wö�c�_�u'Q$��f#Y��U/%��߉ FiD(��fT�2Zy�'ҝU����@8#�]��v�R�ɾ���78@HZZ�$�e�����=��;4/	�L�bM;HW7Vêp����J�eo����o�j��D���q{�6rS����0�g�	 `� ���g���.���ʡϺ��̾�����U�3�YQ�l	�[��$��^����.~�������H���p#���:����Ҫ��:��:�G�� �t�,���E�5^��9��ܢt�	�mǛl �Pw�(�*C�hE{5P�&2�\_ŎA7E<O]�A�S��ŧik���<��pb�QpӤ�Y,k����'C%
ttEg�-��D�Ɋ
8���(��{�����}�[f"5`n��~܄b��B��G�a|4Q���R��^M�fxV\��g4eg\1�x��`2�����:W��t����C�d��I��Ma��:1����	\�G����{ R�~pPS�X:B��Ux0�0`۴�~��v"�\r�9��̫�y/A��̚"���0?�h�aw3�x=*X��L���h�je�xO�;�v� ��,��o�h��̇��SĴH�bYm�!@C����~�&Z���J{�,��$�D�Ӭ'�@q4��o��11��di)��p��fN�/���.'N̘x���"�m��a�F �5M�,��S�V'�u�F+k��Ý��A&n P�p��_���w�ɩ���1����X�Є�ǟ�d �ç{�O�&T]��m.ڈ��'A���oF��|Ά��8k$�a�c�w�"�Q��_�Ija�P�H���_�N�NH~�<��E�泝��!����<Yb�!�H/YN$�x��l �Lc�!4`:q�蠥�G��m߂6�Hmd�_+�T�/��>�LT�zH�
�c��qC�,l�7i���o�+���䧭��H�����^�/�*�����z0Y��0�Ǹ7#��O8�bف�dm�Q�`����9&Y����
l	��y�n(���G�I�x7��$��0�^8^�%�H;J߃BD�I4q�T�T�����ß3��#bl>�r\pgZf�'Eg���8�̬��N�x�����%)����� ކ�����V4Y�<S�Cǽ�T����}v08�E��:x$ +~�u%;�����vwPd9b`b/�ehn�L�*�����1�F
>��Mf�?�H��G,}��:r��o!/pZA+�m.��,��O�H3���)< 3c��ܫ��I�`������OSD:��T�^emz@ڥ;~�t��� =��� ��b!�h��ddL�Rc��A���썰YW%e\^����k& ��h�R@�MJ�~���g?x�(�;��1��?��\�d�z��a�ӂ^h�-nH�*���D�Q������G�4��O���g��{6�j�S��煔�x�v�Ő�$v�����Q5v��iu��A[�T�#��ߒb���`�ak����rM�ҿ�W���/p��N�/��_�>pE� x��H����P yE
��/�(_�z�C���/w���F6�8)N4|��gD#�}A#���~�����������S�3���8��Lf���e��2NBk����1&fi�W��:8�XW���+����X�Ő��4���:����@!|��<0'�Cvٯ�ЊiGLylg�ND}1��,Uv ����#̂��1t�T	��ժ-Џ�v�nf�H1�۲��SXZ#�Q�G�.IV�W���?=Jk�_8|<u�^⯿��]�if���1���]k��v\��+#�(���W�T�:�&�>�$46���0���Pd��eR��YG�+�@�����ʈ���(Zˬ�@���F�,��4��>�[]}#�˥�X���XV��:+���J�h����d-H�$8#��n�%^.��`;�8�fYj��N�;|��@q+
��n"��ˣ� 3�~��Y�	(�=@���!��߁�0��ia�N�vƲ�cZz��i<�,5Cux�>��d�s酑�7�'v���
m�bY'
��wl���Z1��1DSo��܊Ҷ.	$۱�I��_ QQ�PH`�
YHݏO�=��em���f
����g��=n�����a��r����V�C�7�IH�L���B�5��I���q�ުȇ*�٨��AL�����bp{���p����u�~ҁ�"���y(�����=j}Su	>��l"!1�%ܚ�z͍��J��3�D����k���g� A|��;����Q���[~ּ�����Ƨ}�<���'�V)�N�=�����$�!
��*Y��h�K��xL�1�Ҧ�E���)��/z�0;��>C/�	�|P�ѡȯm����������i���
o`'$Ț�z����}i�(�n�SU_�k��mFK�U�?�qyO|��	�θN�;m]ٺp@�I�&��1H�"�e�$E��pyo��0�l�<��$o�t��Z}�"�sxll�h�Y�S�]S�J����{`�ܧ�D�5-U��i�
]v��?���z������T]��v̀pF�C���t��wΆW��t�	]�D'��N��cE�It荁�Ǐ�����?�TuL� �eyCx�m��|�}5�UB��,����{n�� �ё��Ŧ܏\P�Szۋ/�}g\ ��{���v��q1�痑�9�<K'�B1��PA�ț�U؊�>�����8#ܙ8>�Ĩط��i�x0�R���L\��xV����b�ޱ��_ɺb�*06s�VBym9�D�U�3�����,�f#��b7��`HM��M6��ؚW]$e�X=���d�֥�e���{]��*s�㌡�.*p;!�V��T(f��}�oht��NH�Z�[zF��h��`/����Q�M�Z���Nޫݡ��%�.���C�o�z![�=k�I���/��A�����p�������r�bF�%�me�PD�2݄K��c��bY��m]��(��o�] Js����*�E����V�p�V@Q}9JҎ���мǰ�XV �Ŵ�!����M�tsW2�q�����1L?%-?�ӡWl2�%y�5�e��îĲF
�1!:�%������~�x}����Ʀ�TO*�ǲM⭶�=��-�s<N�����x1?�k�O�J�`eCTwqE�wG[��je�9�gL�,�G�}� �ń��0yYdT����J�(��vJW���)	�êW�@o]V�\۷�,�"�(Ꮁ��:<.�i�/:�"wn���2�]��5��~yBE<h2�TM�E���� (IZ���ȃ�8�_^�&pLq(����O{-Cл����-���
_oZ��^�k]�5A:~�!!=x?J7�g���T�C5>���^g�@SԕVAx���x���v�Cbpe���o&?o`���_3��qz�!e_ğ_;�!��3�X��!���A9�!�pN�(nJT�0���W��;����Q<�d��L$�b�-�:�&�ĳ�����-��$:�=��q�yhr���[V$��2P��=��ux�c�����3囘Q�L���z���K�H4�h�7�)�c�Y䎦$t��.͟��6׮(��K��� ��p�ԋ`O�!��4d���nJ�f��I�A�5��`���?.�%�	�q0��S��M��jf���8��E�E�n�4��-�qf��u^ϣb<�Sq�V�Xy�!3/�O��$���PW�FX���,6��NL�����v
�hl|��J�84$!
�-��{ =��I�%��8�e*8�� �n4�O�o^uO�,�ucb����u�@�UPS��y�n��O�{�W|UŝceqTs�֪>p�gk�ef~ʋpny�����|P �! �unU�WU�Y�s�m�Z'���	4W��_'K���,$@qm9S�Rs��n����m.�&@��CT��p@��:��b�z,����xg�[����(��.�M���yYZ ds����~G9�ǲ�6�-ܱ��QD���?�*���'����wë��>�v��&_[���[~��+�kf�S()�5�$�5���E@���\*�)PJ���'7	2&�?\8|
�e/�� ��R`���p9���.͆��� �!�q�Ɏ�æ��n�,�g�UH��E"ю���h�~XU����T�Gl+P�d�k
�Qe W���a��A/�#���SxU?�#�be�_�s@CgP��z�p��zhG��FQI�<b������>Ǭ�&Xl�
���xQ���u����̔ܤ��Ԟ��G=����6ն}�"p�bg�Z|h�E��w�A :r���,D�,�豖��J�{}�ϻ+Y2\g�炧�KUT����ﯓ}��LtXض6����?�;���A,s�ʜafۋF}{���~�=��������ܺ!����'�Т����tở��R��y��?9���cg�o�9��)t�h`��|f�pa
�;��h�������U�:�լ+���(��
�l>hӧ��[�P�[U?t��$�x�����	׈�>(o�2�?޸$b���F�ͣN���Z����G�}�A8���)�	T��=��]?7T_g�)�{�1��b������;Q�C�$��sQ��()���zXH{�[edk������0u��Qt v��l	�ŦO�:���	ҽ�e;��.�-�Q�J}Y� 2��JQ.�X����^���BVT����b&
e[d�E�B�A�?'f��%�U���g2�eƺ��緟:d�J�+��c����,�7V��",��\�����/�^/���T|�DVNe!�}ʥM{-���/���ep�����1}8*Kt厈�V��w�e���v�&c�_
���UT�~G(��e1����
U�Xϡ�ށ�!rޠ��ࢿ���"օzcU@w�g8�u�����	�D�؁���:��"KL��,��pƑC;�1�=���ڬ����f𼨘�h��u^��a2���A��8r�	��`����&m:�E��\}��>a�t Y�2{?�.iUH�	T��f��'7W$��k�*$��LnQME�Q��#|���3�W�V�_��<�&��'��_��J�7H�V�	q��Y�E;�B%mC�tңU��S�Z�d�a�<�[5=���Ǡ]�����D��8/>&��j�U��}Jrx�o�����z=�J��je�����<a��4��[Sz?��C���ߩ*��-ѳ�G�Ց=hM���l&<|�5,����5/�ȹ��@�xʊ�D�����S���˫.����M���N�[�����G�Bϸ$���i�,�2��[z<�rK��cH#�c�q����r`��L�|�Ͳ�i�g�'*h.��mfA��B��T�i���/94��6����;f�	�c*�� ��Tӟ�τi��uZ��(>4،0k�Y0��V-	JY-��@'�Q�[�u����/���?5F������#&�3��=c� ۠:±�(V�(�de�]wp˖�r�r�R��cT��14Lh��k������.��n�]FN�N-��G� >�����rn�vGí���(^���/�P��-�H�1�d�	�q1(�	=�����{�>�i��p練� t,7!�}����
��.aiF"�GU�N8�:�x��[�ʹ����M���{�������݋w��ow��E9,_��{g+����X���.��:�*x�w��O�߆p��IQ���q�	q�����*�S�P�h�(=�o�?,��l$@h��`�7O��=���v٥��e��6�!Kwo���W��Y�C�����ęC1,�/\���a��_�9���!���T�	a{�nX���WR:\q�L�����W������`5���w�ow���n�
4�6�ǖ
��/"�=w�mp���t��XVM$��L��I�!l��$�����@\�����*d'!��e%S~�>���)�M@��ଫ�{��w�#���JL��{1�&&��S��S��;�3�^~M)<��[o��Gϼ�8)Qo�?������Đ_�(�b�6h�K��������"�z�.�Q������ S�+JɁm-���{�ĝ���j���
!�k���q���u�h�������S�DPM�C��GLLp^�A������B��h��+�}.{*���[؋���	fT�'�f|n[�~��Q�h��Oš�5=?�й��(P����EU�E4�^��~v�m�}g�B(�)k�
��t�1��8"��N���^9��PP]g?	�5�N�q�F�	E$�*�&��M:l�_1�E+�K&�c��������[ݨ_���J� 4���B��,�X��]�Qd�i�Mۢ�(`�m|�ۏ���o��Ɯ�/����!E�m�,�-��w��_�2�Txb��PB�؀�ݰ)j�=2s8<r浰%?�^<\�F���D�a���oROx�w�&X�j#��+�z��ꩶmྦ#W�	x!�k�i=��;^���5je|����z.>�,�������A��
�>�5��̫�h7�M�΃��֓qA".��F��������/p�ⱆ�Ų�Dz
�v��SZ��À��k�p�
S[���鄀#��k�K?`�q��(�~��T�7Q�7~��e1K5Z|ǋ��	��^`��þ�8��������[]獚
z�h����c��>�a����R���VN/��F.�/����U�)�ߠ��������̾_���- ���)GxL����Gn��Yx�����7��z�>(�*		��}���i2{�(��a��j&>?k����'��o�����cLʝ�M'"�$�|��-�i�(�U�O�n<�;����vU��{zLҿ\���uhc��<߫N8Sw^��ˎ����[32�PW\��n���̤���[ĩH������M�r(L�7
������18���R�q:������>>��
�}N\
 ߃u�o:�7y��`Lz4uc���8��e�k'I�-��"�OS7�w�ӷ>��#`�ߜ��2��ďu��#�������&E�-G�2��~��
�Ε����o��sJ(E��	��J���`e�K�I�^q��w���+�m��h�����&���'.��s&Ύq���⍷�P,k��m��|����ʜ{�#���{К� n����ê;N#�=A�Cj�{��[�#�JED�1[D���Mb��k'~���A4g	���>p�uЈ&6�NY�/����ؤOȡ���'!w�E�V#*�I�`h�>����Y�����;rã�@8#�a��������;L2h�n�^II�b��Dſc�b�E����j������{H�t����u��d)���g\͂u��A��WC~UO���>	��:u���(�J(��zcԠq��}��,�ٸ��)[�h�%[W2_�˛�a�5���Y�Ҋ�!U��}�����o=K��|̫N����(a�.��W�\���l0P��i�{���*�&������i!h6E��7��y��`�y\�����߈�=��ٛ�b41�:�W�/�)�m��� d1���|�v��4X:xo}rPD}CIy���T#C���,|�?9���p�(N��Ь^�J|!���Q�����,��$M�z͛�8:lL��Uw�QUY��6%eR 	-���J"MA,A�uU,6\�Uq�UV��(*� @�D齇:$B��$S��?�̈́I2i����7�y��{��s�i�E�ۍI��}���}{Kڲ�ѤƕI��e�A���Bh��sre�-�l6g��L�YكXڲ~
-2�=lR��u��"屨����FW��c��S�%���Mq���F�~��<��H�ɋ���5�������Nm���xU���˗��Oqzj!ނ�9Y�ز��-O�h����6�O��P���TUW�)"��_mxX~��G�:����z�H�`�|�����y7�`�X�רEC;�*b�ϰ��{��l2e瞣L�/6.��!�ڠ �LBW����6۳��cز\���lY�b�˻��.�~Y�=p-[j�pz۶�?<���;�&�,ݻ�H�`��cFCjz����S��WX ��\,y�����Ohج�h�����#=��yl��o��oN���`�������#����\��v7Ш��ҍ-:�|�#?�L��Hdo����Z2�o��\����C�/�< z˴��AZ��w�����{�#���S�a�W���[��rmYR�?�VvBL�V*3��Wg�Yd���,R��ѫ�Ǌ��!����sb��Ӟ�M6�$pi��h�WSh���L.߇�WL��g~s����E/�]�����A���f�"��2=I5�H��$9I3K�09�_�]��Ƴ��F���d�u�U�-p��Z@fx���H����q1}<�9�`��Ȉ(�[ �I������"�A���aV��J?n_E����_xn����̓�
��xg,]-�Uݍ��Xl�*'Y}�z�f�P�&�N��y3#vx�T�%��M�vR}Q�ck�qFp�?���En�@Ə��Р�I�e�K���l�LG	��	��I0BX�/�9̯�,a熭�Wnu��Z��7��+=�x%`�I��x��Zd�(�G���5h�����3IR�����rQ�Y�00��^]����W�>-�AC��J.����J!�/	J%�*6}<5�=�򊝕@�2��,�	dF΍k)��N�9�uR�O��<��:	��?q�&GY�N~8��H�j8��W�~�6���2K�ݡ�ܺ�J�k\����jj�����1ݿk��MC�yU�}]T��Uy�E2.� p��s�`��0�����k�={�0ib���o���3�r�ׁ�D���uk5ۮ�2)�t�b0���b�����u�0J=S����s�`�.�����V�ۢ}KM��5��s��%+�T'��_׏�:/�;�y��-�9'R�)�t�sĳM�S2���D��[���%�%$�[^�� +l(L�����n���7>��q1��2[K��
#��D��ш���<���sWwh���\���0#��(߶��;�.<����y�?��}�E{�2%*~<T��|G*I=8��#9e�g��mf�|�=OJƩ���X�\�u(�I�T����U�7�"�A�$HN$H	��kt�K�}?��(F.	w ��c�=���/�M u{�w���8��jԥ'n�G|��v#Z��>(:�Y�y�IS�ƅ�N�<^aw���0=�ٹ\z�ȖŰ��?a�O���1��TI*^���$��>�Ȩ��q%.೐p� ��.w���l"������C;*�� ��L����oA
$!�C���РF-q����Z�{�/|<c��?F����7+pS�6�����c��p�pie%���mޞ�=����q��.�-���[�k\��ڙ�n�e�������D�tU���&U{n�m�;�����\�H�6��d�ڕ[�;Гy����t0��p
^$�P�*�_��¥3���5����ia�wtw��EZ��@����Ә�w���nM�|��ş؞P�M )���A������7��i�P���b��nk݅%5���Oӄ[F��@n�+���魳�\�;���%�Q��/x���^�s�Y�e�ʋ�*�/p�'�9��&aob͚�&�۲��	���i�ϟ�g��HS�<I)��_!u���d$2�xW2ۨ���0m`��b~A>=�՛�N�[G�r��ƻ����;�KT�=�%�`ϥ��5]�S�:T���ǢY��R�j:y�_��e�Ю��	�2cn�ʬ6H;��]$<MXJb�y����a�@����(r=����k	�,�5�v(��	"�{��>u�x=n=q����%6���>['T[�PةF[�(l�ΐs��^٢`�ٷ���{�g	�,���8�~ڳ��y�R����z`k��Rr�w6�'¤�ϴ�s�H�;r��ۦ-޻.P���o�ڲ*�V�t 0���HiǄ�K/�~��r��,�����Z�K�r����:T�{,�n�`<�~�?B��V&!e�X	�.��P��q�m�)�3�_�u��ٖ	N�h�=*��:�]��x�r�o><bG5�����+��CC������q�g�tbi��#�$H�\]b>�Z�;�l�~W�]���]%�v1 ���r#�e��I- �&��ޣ���:M��0(��%L�mH
�0��>쎉�G�Gk�C"ô]U�G'!7��Lk�q2�> �=$*��!OO]@�g��w����p�{�vL�l�ϥ5vX,�1�'{m�gW�pJ��'k5&,z
���ؖ�Q�$?	�����l"Y����P$��UQ��I#+&�#:���!1EY"�NRei�h.4�nEv�OSWͣ�S|{�C�X��P�8dH�^N��/x��p�=Hl������{�-����]��?BV<��o�G�o3I�pM�z��\?RH�s��i�^ώ��79pld�-�ɼ�F[͂XU�
�C�T�(���y����y��SBUW�z>eٗ�\��i��!=G���Kq��k��`º�'���*vk٬ݳbȉp��6�I'���C����A�c��v^Uϓ�܉�I�%�hu�4쒧��~��Z�'.q�&Q��>��~���U���O��2�s�8�!��Q��s�NSϘ�l��!�]��,����'0��*�̀�3	RU�uDhB*�8�u�}: )c�� ���v�a�dR���R<Ɵ�`�'�,N�7FT#]�u�e!#�M���Ę�^8��ev�����s��ZH$�+8�q��jJ�n.��<�m����֞7F
 ��BR��NG�a	�֬�=�:"�A1�po�C��ԏ��k�+��"�))���\մ@ '#�A6�?�������b�;�#l�U��++KS���3*؄�����l��ټ�������o�N�8Z<k\���]Ǌ�q�[���X|!`:Ph_44�^.���hE��p/dm�cMR��K���T��\ܖe3��%����#c⥍؅4��/Q�%�~ؽF8��:N��h���tY�� @p���}q8���GāR��E]�f���O.�~��aJݵ����m{n�`���6e����9t�s]V� �а�Us��^S�sD$��R���#b���ji�N�w�D����1���A�A��c�3_��^¾HQ��3�c'��0�%{׃A�ō�wSD��? ׋t�f:QwЇ�Ј.��]��jnL�
y�/�و'���-�����M��{�
��z+b\��svc!\KP~��2e'I�l��"3u���!5���1��B_'N`�L;JìXi�-�g��#?X��!�TW���Y�l��y]_q��<������8:7�CD�&���}6�sH5{��m��n��n�n ava��(��x���J��0*jl��^n����`0n/2�f��em�:���9��.�T�����@N�6�i���!e�<����u�E8Zs-��߾k(}�#�+�ar�����f���pS�,�Aͺ4
$e�+[f\}=M^�	+��x�^����Np��������M��7�^\���n��-�C2ީW*��
e��,��,��܆߰�S�T�g��}����+�N �i}檹�Ъ1�@؍��/���y�CԪ��$�	��*�R)I:��H�]��Y �����Ǚ3p�hCA��1\U��PH�$q�&TQ\w��a1���SI�G�X=l�*���}�Z���x7
E�tl�q0տ�2L����T������T_���ZU2F����vqO[Q-�R����1��E��K�6V���!���y� !|�ZۍJH	�YZ��4C���(�n�L	R���o��?�6�E���	�t��ςV��,�����%ty�ޙB�o#d2�����ࡺG׏�v��i�[�9���+��M��ґ��V��X���x83A5�=�.����m"m[�06�>�=����ޗ�\���7�:�q�F=��ؚ�C�������EZ�DA�g�"�^AfƗ/$�I�\�ï2Z0�M�P��WБ"(���{��rU�+ل�#QQ�~�RѼt2�lv\�i�i ���iN���Y^W~D�E,����4[��5T
 ��BR��kf����̣��;�qm��7z�b��tU��j�/��Qh_�u@6d�*��WW<h/���c�\QDA{޴cryN;�F������&"xJ����@Y��@َ\���X��S<��VI^j�A@Dg�eڛ�Rn�l &�,	�ea�M-�ff��7���
�mAy�\�E�Y��u�m����-�S����,M��:&�
����ᤆ��>_�r2��1�x�������Rr�,��"�DiY*}��J37Y��ʰ�ܶ�[��*�����{��(�W!m=�F�}�D5���o�7ӈ����?�]n��{�������1�\_u`K��3쏣�uҸk�e��4͘���$�W;��������/��-�Ilx�:� �� �����n���	�s�z��9��,��`�	���l���@�:S��d�M�����RJ������5�����:�>�C}S\4|����劑"<"�"��J ��>P�c�>�l�bɎݍ�Q��;D �X��-������x��Jջ2�˿�G}Z��w?HVp^�q>z�f�q����:�v��J#0;R࠷3ҩ[t\�x�Ԧ[�*�}7�?y��}Y'���)<=	I fЍ�jݟC�k���6�0B@���`{[�n�}yb�(y�����B���ΚѱtMrs�Ȁ�@��v��fd�^����U�Bg�׍�%
���n�)��#�GlE�|Y����o2��ͽyء.1/�Ҽ8�܏yE��Rj0�1#���WJ/6���<QԠ��꺛�^>1���a9ǭ�o�S�����pKks�72�����5#�1���7�><�'�Л+"A��� ��@�i�PW8O|�aиƮ=����V\��sv#b����TA���Iv�L{����-��9:�Q���E��V蕎�J�f;�T��M�򷎵�#4��d�a��4;&�3+L�ùߥ?`����M�1h��x��%���=۠M��y#��L�#���Le�UI�UVUoʿ�<<%���]�~�b&}�q����%0j��Qd�14������2�a!J���;��?��P
]bA�x�<V^�W:�7S镒�;��\H�M?vݴإk��|e��3�rQ��,���/��A3V��a��n�&��U��Q^z�2~�|��i�	3��^��c!5��I�������L�������4sٕa��U/�\ѳ���L!�˳R]�Z��`�,TrqQ{�x�I[�����Գ��~��=vQ�"��SS(�aѻ��65]F������E�����,�����R$Y�O�ڮ�#��uѴ��w�)�\Ւ�������f�~NQ��K0	Z�/ܸ���F*�Z2���3��"�ԈK-���.�в��0v�o< ���(�Z%���:{z^�y�AO�m+�IXVl J'��dݭY�����
����ٖ�Kx"�%d��9ؑ
dȸt|;��4ڸ��ȑ]��P!��XԒ.���H� )q��͎Z�w�s�k�>�b)��������E���9�1	�12VToއ>Ks�N
R�Cļ_���:�#�A����m��4�W�QPs7Z�xS�r0�F=m5E2��XK�M����)��X�<���솺���fn��y���NҶ�4~��&����6Ӱ�.w���ԣ�Aq}GZS�1C5�ɚ�'�m�Y_HH�v1�P�f㮭����H�|*X���X����q����U�,�4IrL*��J�` ���$ �����#��If�T}S
�- s���zV��'�rM����oۚA,���o�M�z4��l�\�xo��Xz0Aĥ,t����JHL�d�;ۭ��TM$=~��^���7O�:on`�f6�����ٷ�$߁]*��=�Ѹ���1�	7�����=�E&�!����}V�rt^R �}�)� �A�@,mc�y3=�{ ��l���yvw��� "��|=��.��mS��|��WM�J�xbo�Lݣ���OG+�tN���q-�;���F�i�\���Ӫ#�bsR�||���LxT�.Xi�	��������1��7�=^\h`1��J��kԈ]Prڧ7�Dn�&�X�t��~��jZ���r>u=/`85�������b2���Loo��c���p&)Π+)��%�t��
�zF�H����uC��s(�ĮhJM׬um��!"�h}	�\�f���j��) <�n��nhe/���C���
��4�gt���yS9t�'�՗���p�F%�AX��>����<��˱��-�l�fNN������2TZyX���Bz�6�cΝU�V�^k�l-0�(�!:}��P����C ��K�A�c�PM����57Ӝ}�e��!�!�ׯ�>�9���p3��Ad���y����k?��,�>�A���b�,��llϗWFҧCr��VSdb��K{V��
��������bR�f���؝2������ϫ�9*涚�ia���)O�]T���O1��60I3}Ŀ���-\V���"˃뙬��7���mxgr)���MZE74�DZ!Q�E�/������|y-$/��ո-�ڙ�!yH��Э.2�*ү[G�54��{z��Kg<�f�4s��؛y@=�u�����XU��-�RR�ٲ��:��ѭ@º���Yږ���hRɄ��k(���V�:^&�� �l�� ���.��P�g.���}�E�/*BV���J��(�_�z��������������nWgӎw0��K)�b�<�χ�	���.HX30�f��%�����Y�-��]��a76����<�W�%�,�b�&��+^1}���ܮf��!�ƖUj���IG�|��b@��c�
�t��j�������q�sZ��?E�\���Ѕ�$IQVI��r牴���dc+�Y���3l���b�s���k�6u=��2.*�2vƇ���1z/�(�����h]˰eYe�����*ܗqL��>�LSV��a[``������i�n��n����
-=h������5�� ��~�е���{��z�!�K�e�	���F%�ǔ�t�u�~3]��ү�K(}��/yW�ɕ)
��=f:���o�ұ��Ţ.c>��~Y>�L��tX^�OE�A�2rd��j�i�Y��0*��(��o�LX7�������"��i�U�{I��-Vј���r(���!]�����.�� �V=Ĥ�����T +��a&YX��h�4��O��y8�[��b��[-������/r���A���r���fL�f侊����˕�����_�[�������?�N�5[��L����d� ��)��!Y���%���I�]�'Dk�)�|��5����� ��vW����櫥+v��Y�#��n���؁�����*�mY�yU������!��mO��    IEND�B`�PK
     Y�#\1�9�c  c  /   images/c3d75dd9-81e0-4ecb-9109-310dbcf70c9d.png�PNG

   IHDR       ��S:   �PLTE�����鼽������껽������������߿����������������������������ȹ����������ݽ�������������������������������������������������������������������������������������������������������������츺������f�   	pHYs  �  ��+  !iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 5.5-c014 79.151481, 2013/03/13-12:09:15        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stRef="http://ns.adobe.com/xap/1.0/sType/ResourceRef#" xmp:CreatorTool="Adobe Photoshop CC (Windows)" xmpMM:InstanceID="xmp.iid:0AAAC2C94DA211E49B7DDEC391758443" xmpMM:DocumentID="xmp.did:0AAAC2CA4DA211E49B7DDEC391758443"> <xmpMM:DerivedFrom stRef:instanceID="xmp.iid:0AAAC2C74DA211E49B7DDEC391758443" stRef:documentID="xmp.did:0AAAC2C84DA211E49B7DDEC391758443"/> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>r+�   tEXtSoftware Adobe ImageReadyq�e<  �IDATx���͎�8�� E^H%��{T����/m��n�HBb����74�<c��npQ                                                                                                                  @8��_��K��nW������~�I���]}�/�?���j#�]j^?�� �����O-������G��O,m����r��sJ���i��cm��)��[i�<^��:�m|�\����ѣ�S/��ɤC�4�<�t\�弃��V˞�g�Y�4�v@�:>xC�X����Dڿ��4��4����8�q0t���ep�mO`��q:�8:x��b�v�@|���'�:�/��!�v�w�U�7�ɑ�8���q��qx����ǝqx����:w��g ���8>�At�+�W8�+���#D�>\q����l\�\���9��w�I�S��w������#<��ZX�
.JV<�+��W�Kn�u�Fڼ۟.J�!;;�Y�'2`beQ�L��d����ه.;��uxǉ�t�<+w���J����G��\�"�7���p}�hOS�Fĕ^�����K{a�8����ְ���j���ۯb�f{X.���,cyܦ[m�>�È�,m֧��������۲�m�\����$���z������{�i����Տ����pܿ6�����J���j�l�t���������+���R����%��lfE����h��)��so���:k�������"��K��_m|.�3ً����ơ�M���a���n��m;��?��I>�{�jsa�S���Pu������c�A|�uP�+�7��׬ҕ�=&�T�\��l�A����Su���_�r������[�����/������;m��ٻ�lBێ9��A�n/GՎzP0��M�b����vF��|!���10[KQ�޻���wu0W����v�f(eo���3G�s��ǭ:�O�q��{�]u40+[�N������AE��ةƍ>ߥ椻�����\t�S_a-9N��^��7���Ƶ}˙��#5�}��8�O��*�'��T1���1n|}�aa�`��,`������z�s�]uXd�G�z�#��o6�(�m�~7���L=����rc����j�w�3����EM�����:(o6k�t��e�@JK۷y��5v��AQ3j�k�X���:�(�'����uP��\����Ľ���?��r
:�o*��L��n��,�@1����@               R�����(��?uI�EK/�5I��E�Kq�Eň�6�(F�G1⨍8�Gm�Q�8j#�b�Qq#�ڈ�q�Fň�6�(F�G1⨍8�Gm�Q�8j#�b�Qq#�ڈ�q�Fň�6�(F�G1⨍8�Gm�Q�8j#�b�Qq#�ڈ�q�Fň�6�(F�G1⨍8�Gm�Q�8j#�b�Qq#�ڈ�q�Fň�6�(F�G1⨍8�Gm���r�8b���m�e�∩o��v�Eͪ��!���c�I��Wq�4 �����8FGT�MQ�c4qD%����8FGT�MQ�c4qD%����8FGT�MQ�c4qD%����8FGT�MQ�c4qD%����8FGT�MQ�#��D#����qJb���W��~��4�
GT%�H�������
h˷�a��CQe�#��a�<[�+��af�GT��8���w���>Ny4!�#��q��g�?�G�ɕ8��Gz]�Xe�mׯ�GT9�H���æ]�!��r�qx�:j�š��8��ǡ��m[�*[��kS� u�#�\q���!�����CQe�#���;b>��}�u�#�Lql����iT���#�<q�N8�����qD�%���ǲꛁ�*OC�8}�N�O�8�����l�z�#�q;������:�U�8�\������*Ci��bU��!��r�1xV�9�j�%��2ıY�G�+��#�ql�w�Q��*qD5}}��o�_�}@qD�!��]q��Z�#�q�3rqD��� q�9�Bg1�*ni[�XGTq�hօ.�#��W�ұm?�L��U�8�w�1���[zbKQe�c���}��S��gXʼ�.��r<[�~��#?�����"#��s|��.ϯz)�T�8��������IW�N��}l��O��U�8^?�;��#Ʈ+qD����/t��I���_���(����1�NG;�5���%�[��8�ʳ����cځ�۷g�X�#�<��:�8��}�}=EqD�i!�ACǤǿ�&�.|�8bʴ���V���}���7g�X�#�\�s��1��5���<�GTٶ=��޼f�I����N��U�8��^վm'����e��N��U�3���?���k�N��Uƭ��o��ɞژ���}c��U�8>gV��v�c6�Xk1��JQ匣i7w�i��iW�q��.���GTy�H���iؘ���۫��b%����q���B���<n�mc��㴯���8����6���>>�XO�F�ձl+qD�=���c�����a?�r���e�X�#�q��$m����n�^����&M���wt_7�3�GTE����5��gǜL+qDU,��z=��gb%��bđ~�<>sL��U�8z�>�e�AqD"�����X�#�q����0�GT�H�E�X�#� q��|���8�
�nH�X�#�������+qDU{i;|��8�c�q�����E�S�&��fG:�]!ݳu�ķ����|����ؑ^_�c1�6��j�q|��׮������SO��������ԩ����I���t�_#��f���]�븼�g��3��JQ�.�?v�1�*��&V�jvq�]��c=��	�X�#����׶L7�����g�4���j^q|��TǵC8��T�L�ͬ8��U�����]�����X���"qD5�8��������g=��JQ�(��o�_�Y����8&�X�#���q�$���q��o�<��JQ�&���v�~��L��T+qD5�8n�`�s٫�揚db%��fǍ���V�諸>y���8��I��ձ���i&V�jqt���k��*��`�YqD5�8��8���ڟ�~�8��C���ul��1��JQ� �~�����zSSN�����X�#�ı}�up�/�uZ���/��GT����4鳎��}�ȉ�8�z|�O!>��M���+V���q9�h��E#'V���q�ݯ��?�����ǎ�X�#���1b��)��X�#���q��5�GT��#ǥ�;�?�:���Q�\qD��8��ρ�3bb%��8r̩�1W�����8̪�K �#�Gő��b%���Lnp�k��fVQ=&���mf��C��e���9�GT��cN78�r��JQ= ������X�#�ıYϴ�;'V��q|̶��ϼc74qDU<�t�qwM��U�8�ݟf^n�s�'�#��q��ǹv�6�∪li��w�<c%����1������CQ��#M�S~'V∪`i�78��b%��J�U�1���8�*Ǽop�m��JQ�c~o7]7슕8�*��op�e��∪P��87�V�8�*�L�n��]���∪Hi�^W�&V∪�ȱ���!+qDU"�M}m�~���g∪D]�=�{b%����Q�Ϳs�˾_�*{s�����OGT����4w�9�GT���ǹ�+qD�7�*�n����JQe�#m�5��sb%�����q:�{L��U�8>*o��V`���*c����K���8��G���tDw�!����Q��M�u�pqD�+���n��sb%��2�Q��s�+qD�'�
�n��]77�GTy�ج㴱h;&V�*O���X�#�,qB�ѵ�8��G�����6��*C�6¹u\�#������o�+GP9�U!�����[-G#���1�8��h�J��#*q�&���1�8��h�J��#*q�&���1�8��h�J��#*q�&���1�8��h�J��#*q�&���1�8��h�J��#*q�&���1�8��h�J��#��q]�m��w�W�S�8-W��7(��􎃱�Qq#�ڈ�q�Fň�6�(F�G1⨍8�Gm�Q�8j#�b�Qq#�ڈ�q�Fň�6�(F�G1⨍8�Gm�Q�8j#�b�Qq#�ڈ�q�Fň�6�(F�G1⨍8�Gm�Q�8j#�b�Qq#�ڈ�q�Fň�6�(F�G1⨍8�Gm�Q�8j#�b�Qq#�ڈ�q�Fň�6�(F�I+�Ė�"���ՒR�U�l)�                                                                                                                                                                                              �����ѿ{�    IEND�B`�PK
     Y�#\�Q��"  "  /   images/c7f8a6b2-5f4f-47a7-84b3-7bbc451b7ab1.png�PNG

   IHDR   d   d   G<ef   �PLTE�����鼽������껽������������߿����������������������������ȹ����������ݽ�������������������������������������������������������������������������������������������������������������츺������f�   	pHYs  �  ��+  !iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 5.5-c014 79.151481, 2013/03/13-12:09:15        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stRef="http://ns.adobe.com/xap/1.0/sType/ResourceRef#" xmp:CreatorTool="Adobe Photoshop CC (Windows)" xmpMM:InstanceID="xmp.iid:0AAAC2C94DA211E49B7DDEC391758443" xmpMM:DocumentID="xmp.did:0AAAC2CA4DA211E49B7DDEC391758443"> <xmpMM:DerivedFrom stRef:instanceID="xmp.iid:0AAAC2C74DA211E49B7DDEC391758443" stRef:documentID="xmp.did:0AAAC2C84DA211E49B7DDEC391758443"/> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>r+�   tEXtSoftware Adobe ImageReadyq�e<  �IDATx�혽��0�a��K$�,�{����K �p�W~�N�'�����c�� � g c r+�V�-��� ��?J�O�e��0&e�lP��t�[/39,y�
�����B3e�e�AE�ڤwsX�c���2[b�f�dq����ޛ�/��)X�����[9�p��������o���$�f��dK��J���og%���UtVҏ߅�Z���5ͻ��MR���Y%P���]��%I�P�('�=�K�:!�������5&z1&�b�brI�tD�T��.�H�'	�"�`4�sǷNR�*�P�ܬx%Ph� M�g%u�M�R��*	s*k�[	�@;.�g%Ú[~�	c��-�c��t�։Zq�#ۊ_w�	㒘�v�K��]�!�W�{���ArI����j��]�t�[����=��'�}G���	� � ��|k�Z�:�    IEND�B`�PK
     Y�#\q�,��  �  /   images/be1ff175-690b-4799-aad0-0ab57f9a01ac.png�PNG

   IHDR   �   ^   ��\`   gAMA  ���a   	pHYs  t  t�fx  �IDATx��Q.lK�w�#�H��F�`F�0f�x�N"��w$^��~�dI)��>GU����%��ݻO��U�^U��j��?�Q	хN%��.D�H�"A��.D�H�"A��.D�H�"A��.D�H�"A��.D�H�"A��i	�ctt�����������J��9<<�ggg�����ԢlmmU+++�~Cт<<<T������eU"kkku�����Z__� ���l-I(��X^^��%5ER�pttT��R������XG����Z�&8���[����M����D�(Z���0�$� D����`͋E�[?%Ebmn	P	Tbj�h������q����Pu}}��="�I�(D�T�F� J�*#%T*�Ʌ��������y�^SFu$�7��5��t�q���h��I���۵l�a���b!�,4?D�����=� a�K�@��TH���saa��1���٩+~~��?�8q��(�H4E�RtV%H���	��i:B�\�;�ӗ�;S43D�H�3�14t:�t:����#K��R� �)h:�����{�m<==՟�Ê4�$�xjj*Y�,� \ǚ?����y566V� ��'m�e@�"�"�F��1��������y�8JX�L(f9z}����Z����9l�x��D�0P�6/�L�ŉ2�+g����.H�1�O#,*L�0�"B0��t:�emss3Y��BG��4��Q ��-]��,%�����;��� �}����w�.�NB|e�T�M�w�BXǴ)M�]4�)"�E$��ب�`1h�L��(݂��*�h`KmY�>��aKS�9b$H�E�y!�XSMӣE����"D�	"\$�p� ���.1�^8=���	�Fr��M؎�x��t�&bت���`�ư.�-'�@>���M��`f6�F���E�pѭɟ���z�]�qn�D�^�rntJMvAH��"GWY��"G�rDR"e<s[Y�
�ím'�p�����9��ñ�c�����c9X����\r��7���|����*H<��|^1� �6�XASxp���)A��"hj"97�s+��θ�&�3����l��d�1J����7Z��E�0�-���D599Y���'������)���
)\^GA����xAT/�kۑo�Ro+e���޾U�*2����[�}F��%p�������K��Nn꽾!ߩ��2��-����N6}�׵�q��.|G<��hIT��Q:�\�3;�033��ږ�y����m�ķ��<��?G|�a)�鑒l��%u[�1?�:/� ��o$�g���nI>�?��M���pU�������Na����6Oӆt{<�Ι�@�"�m�e�n�{��@VA����
�t���\��n�!#�47׎YOG�Pp��(4���M�$������
������M��Ʀ�(�m~ƦJ�ce�£�I���5Ʈ����;��7m�f��n�<S߆�b7_c(kw
���D�p3s�)|۪�s�����γ-�5Qf7Z��I��(.�*�B�	"\$�p� �E�	"\$�p� �E�	"\$�p� �E�	"\$�p� �E�	"\$�p� �E�	"\$�p� �E�	"\���{&���    IEND�B`�PK
     Y�#\�Vw�    /   images/a7a20d0b-f771-49dd-a52a-92c84cdc73c6.png�PNG

   IHDR   c   E   ^�X�   gAMA  ���a   	pHYs  t  t�fx  �IDATx���T]Ǐ:v�݁�b�(&����
6bw����b`+�(�(*�������������:��3���E������/����?���?�!#���a�0+�AX1aV��b�� �a�0+�AX1aV��b��ׯ_����r���s�)RDJ�*%Y�f����'��GE�C���Ǐ%Y�d?ׯ_�$G�ҬY3I�2e����ٳ2s�Lٵk���'Oy���|��Y�֭+Æ�-Z$�Z}c�֭ҽ{w�	?�<y��7.�����S-Z$�&M�4i�����B�
�+W.�֭[�Y�6mdԨQ2~���E�]�����B�13��2���v�;wC�J�V�d�ҥ:#��ÇR�L�U���n�Z&N�(S�N��ٳ����úV��H�<��L�.�0@�-*߿��<�,����P���=�Kڸq�dȐA?߻w��$g�e˖MgχT�H���C�f��pfCڴi�K�.R�\���o۶m*F8�p�ʕ���͛�
q���ݻ���2e�dɒE�3F�?.111�jժ��57�(���K��C��.H��r���;�u����v`
��ϯk`Ϟ=U,�U����رca��Z���=y�D�ի�~�l&4=�\7n�3�dɒ���;�ٳg���X�	�,`�CĦ`���*U*�qc��&S�L߽{g����Y�#M�)���XNBPΜ9��ŋ�g?~��ŋ�!T�s�۷O&L����{���9	Y�������kb严`�N�Z�\���?~�(�f͒�y��Mz��X���y�qĉ�=_�|ҤI=�K�������%cƌ:��߿/K�,с��7m���>�����R�D��rO�`�t��I<x���6l� ~��2d���������a���2{�l] �z��m�"0��/_�>�u����Ç�g8x"#�l�o�����'}O	�O�>2g��Au��Y2gάb�;Vsf6�>}Z�.�ڵӁ��Q�fM���S�CX#�4j�������իj_/]�$#F���ŋ˖-[�8�pٲe�
(�e���C�:�F�A�nL�6M�l����ݻw54SA�ر��.��&�3f��~��	uL���y��R�N�8�)\�!@�$�쭗�N+F���{�� <�{��9u���qV+V����)��r�'O���O���)V��ZY�R��L2SJț7o��vO���M�_Ӎ۾}�o���F�5a�Ox"B`�(9�$j������+M�(�E�h۶�ܼy3�q��	�K+V��I�߾}��A�k�ȑ�wps���1���E��o�$p�d΃Ҏ�˗/��i�&��J$��z����,"p@��̴z���q�`�J��o߾Z��ݡC�O���r��֩�ed=�]��^'���Y�F�Ӌ-8�%��i�:B�ST;w��{�����УG-�Pn&k%�-�������{�u�3ᨾ�=:��2���7o��I�71�6@��,�L�`b N+ҽ��\�v�}�N�`P$�"ҫg�X<sSl�G����d�~;Sf�&kF��޽;�/��i�Sb�a8p N���9<���J?�Q���f(3 >��#B��m8�,"��(��nI�l�K���Ή�U�J׮]��B\�s��)�3��aÆک#�ϝ;W�5žw��S:��qܔ��F��M�*�P�f%�jժ鍳���ѣ���]鶱��M�*U���2���-r>'�C��Ҳ����ϓ5������*����]�z���%Zp~?B+3a�ڵ�������x"6uϞ=�\A�E:!���e˖Mr��-���u�x��5�V6 ���{~���bD�6�Ü
�pM�
�P�w^�$q�f�g�� ��-�:I����9x^B�x�Nٲe�e��aV��b�� �a�0+�AX1aV��b�� �a�0+�AX1aV��bĿ~@W�-p�    IEND�B`�PK
     Y�#\�� <   <  /   images/e7e47810-abf9-4bb0-84d9-bf12c3babd78.png�PNG

   IHDR   �   �   ��@8   gAMA  ���a   	pHYs  t  t�fx  ;�IDATx��x\�y%| L�`�w� �{)��
Eɒ,ɒ%Y��I�6�w�X�M�ػ��8�<ٍw�%���Ȗ��E�)��B� ��3�>��MQ1�0 0���5(`���[ϧ

@���

D8�+�x($W�PH� ⡐\A�c�$��|F}}=�^/('bcc�������)?w�$��l8y�4���n_Q�1P� \����ޅM�6B�VO��&ykk~���Q^�M\�:(�+�B�9��%HLL��s?�O�FB�
X�6@�
�{{%T��Y�q|:�G1j����
��$8	7(���
"
�D<�+�x($W�PH� ⡐\A�C!�|@t44�(�Ԁ��'� T($��Q�،����{Q&�>�bA�<Z���$ܓ�Ev�U47���q��-�#��B�:�� �A���~!����N�CCC���������&�l�P�b�1]����P��;<��W/:l>8� RpC�I���vy���cdd.�]]]¢���c��,<�6�����CoI�Jk���7�l�[�@/D*�KrZ���Q����8~�8N�:%�����a�X�i�z���c��[�9��~x�I[Cb����5�ƚ��h�cU����s�����q���e8�(�*�?A���χ>g ޏ�Ę����G����u|� F�~�>z���h�a1Dc�Dx�10DO��}��1�f'��.�F��3�7�����@xk�{�be�ñ "�������ɓ��/���A�r�-���G���'����	�r�Ȉ��M8r�~�ܯ4e#��v��E�F���G��wg"���t=��b�'���ѽ����e�Sz�lږ�۲��ъ�tyl��?v�y�L��%ވ;����f�$�AG�0^y��|
��!�����C�|��;�r��uz=v��ܖ�$yz1<4�߃rO 6���Lعň�cN,^�tk�p�H/����`|��x饗PWW�;v`�ҥHOOGBB�$����j�%3"3S��m���#'q�t:�6!qɝЙ�&|�M�ވ�k�((���_�Tw�X�(���_QP	�W�܄���ۏW�-/Z����f����i��o�cÖ��9Qq��w{ŹҠ�$��Z������L�2҇�E���I&���C�z� ��K���������.��*����T��Ց� u���&`��|8��_�9&�{�Γø�%��
�K6�q�T�y�5ꃸ���>Fr�&~��,�mۆիW###CZ��#I΃ϱę����ç.�T��HZr7��D�L��=,�y�=�FU۟��><��߁���ir�7F�n�kJ4H�G�*�E���*8�o_����� �Z�|�H��`�vQ� �%��6T�{�{�j�.����(NB[��	d��T>���^�<1�
w$I���b4jX�X����v\nv�aD��x��XUv�]�@����� �]�8��@��A�WH��҂ӧO˟w�q6m�$-�tA�&%%	�V8�o���0�[�5��3s^���>0I�9��@S��$�&��!<�Q�
?]��A��A�΋����cn���C{� ��i�	���`O�g�-�y���BoT,�q�|XLш�{p������S�_]����I���V�B�0�}=��k���������!�,\$m ��O��#�p��2G��(:���6lܸ;w7�Lؼi#�"H���.\�$��6X1D��	b
*���2F�iB�j�zj猌2���	R��8)~�^�{d!0�\�Ǌ�
���cѢE���f��b�.**�W��K����@(�E[1��O�$�0�l��^��|-��� F�1H�6Y�7���u�lO;�����7��@P��t,h��I���~���lٲ�J�d&A���;o���qy���v�3���r�͊%�����k��`�bѪv��\�:z��F4���)Od�XbB�m�o��YµwJq��GĲ�6b�"3�]��U����pw�ݱX_��)��.?|��g��I���ڳz�������`գ����X�1�$�R���}�{N
��ln�\�Gi1�������u#��xu�� �6����`]e��F,�� P؊��t�ak�〈��,I�C&/<^q��w�ޣ��������5քۗ���� ��u|�Bݒ��S6$ V�n����؊�"x�r%i�ߣ��0.+M.P<xP*egg��H($�9��ؿߋƲt�_��\A�����n�'N��BY-�>7bTZ������Y�i��\�%��Tk�<��A(�G��<���q����
�����f�-f�ǩ �AL�����c@�4�s�/���4�1�vZz�8X��������@���9Z��h��wxQi�GTh����p��p�F��Ίb��b���?�Ee���AzD��G���GErrrh���ąoF���w߿{~s���ŝ���p6--	�l�����~Sr� �M�x�i���8{����	�t��"�'�1��044�={'Y�5�j����O�೭��&�ۍ�S](��Ku��ى������d�>$�F�)��>����mX|�ԷM-�Ңɟ������6�w\���J�"(PN��Z�SU_��b%j�^n^�[��Ⱦu��jG�`��Eٓ>?)1��²�����*�@�臫T��.��;w�@.JW-�E��z�f���<:,٨X���q7~��ͱ:�]}XEe7Ғ���/j����Q�JJÚ%��R�[��T?Fu�y�jچ�+n��R�#��@��ـ̓����O�IT5Ġ��@~�i�u�;�]=u8w��E`��D��� *zA%)�	PQHr���z�j�N����ڋW��_J*nͫF��Eȥ������ZN)���CŎCN���?q����^�eҷ�=��;�#��?��K�>��8�q?2��'x��!lN����u�B�<�jŊ�w�9�	s��AxΝ�;�X�t9��R���9~�;y�G.�HE/v'&@��>�[Z���5 s�9�@A��bK�K��x��	I>:ԇ��Q��� ��
�>�E�Ȩ���^9��-�P,Z�5�hWw/�"�L�Ϝ{C
"�͛7���_Ggg��B�ހ�7�aU6>��r���,�H_��W9q�L/� s'ג���݃��[���d���'�؅��Ѐ����r-�٫��?��m7x!S�ݸ��u�Ƣ��w�{M@\�J(P0[P����G��'p��a<��c3�&�555�kl�_�	)�P�`��b,����܌cǎ�.�L��|6��g�0Ô�ll�
f	*l���;8 �躰�i��dMM-�|o?.��a*X�e���(�u\);2��YϽ{��>���FQQ������T�L�%A���{Gk`.�zKbT�O�+P0��Xm}Ær#�_��W2�뮻�j�*Itf]�wr#0����n�	���ۨjE�������(%/��&�c�������w�����[��o�����R���LVVք-�>�O
:t/��e�9���܀�M�1Z�+�i��i���<&�M�3+Bѡ��_��l��xG~ �"`������Ām]2�U0��@�=F�he0B������P��i��փ�s�R����Tr�G(s��?�R�)��$ucc�T��K¦.fc�Z�m"�M�7*AU:bM�0%@gJD���>�(|n��qS��sGt�&!���5�GOF�[p�a�Fà����\)Ex�l*++���F���I���D��:ټK�dl����B�S�N��ɳ�k�����%R�Y�_�n����<x����u
2nq9Ŀ�z��eO����h�4Z�5zIxJ�E�tRX�����n_@�#�c ��f)�>$j�a��������x$%����4���-yH	��j=3�Tm�ֺ�������Ty���x�=w	���&,x���T ���v�e��H�E��6�=��d������`�x��f��
z<����Ak����(A�M,�t	�1&@g�@lJTZ�X!u2K%u%�y�O�8H��֣H�����ŭ[�H��#$;eũ����=�܃�۷K/���era �GA澦r�Z��~A�+W�F!�%�1�1��</�BZ� ���&\�غ�e��f����m]h�t
U�4"!�欕��Y�0.�S�O�m�`�~Ļ��{
�V��A���,uM2S���nCuu5~��_���?��8�jQH>M>ػ0�R	{�E8�{Q����K�Qp���HO���F�N'I͋ƃ�=Q�>�,�E,D��+�dy�8�@sk'j�:PW�<>�Sr��	�+D�?4&i�IpG�ص1��}�
db#��T�C��@����������{r��o�]>N!����pO� wt~2�Q�X��8S1��҄uI�;E�s�i�>o��u��ɍ-�=X\�)��.�����6�����,�mB��J�����tQ��~��R��wm��eKCV��4f�Yj�,f�?^����
�C����c\���Z��.��$���%ŋ��I8A�F�3�5�)Jy���FT_�AMmz��0��˚CB��8�ϽK�釽�$JR��o�mX�|ٴ	~5x��-[&���N?�.��;s	T�V�;:Gm�� ,i��a�� m5�^	£��>�#'Π�]q9�R(w����L����ho|�����Gi f��Wc���2��oH������=�ׂ��/ �с5ˋ����J�Tya��P^���w/�lބ�eex���U�Gb��H,��qz��L�.\=7aݚ�X,�i6z��/_.��~�($�\R�Z+`�|��+�ʥ����%ȔpS��D�R�j5?��M��J��K�q����nd��伛>r8�Q��`��7d%\��1+�4F
ɯG_����iÝwoĊe�����ՙI��V�E��H��������? �� Li�r�՛�sH|�X5XRZ2i�ߧ��Ս>�B��J�H�e��."U5��Krqם;���0���_D�Ɲ�p�(.w�c$��>y1��	��yF��`����)�p� )$'8����e넣�0r-^l۴
[�n�|-�;�1/��:.�����AT�
�g�M��߂�8�� <��Ģ�Br��m��m���#�}�jܱc���(R� 9EX���/��;�`��c��iA�ڇe��l! ܥ�xRRB����`씓����]���s���ŗ�kW.��9QQ��	%���8t���-r6�c�-��e�Ve�U��Ă&9{N[+���=�V��kd�2�y۹�%˖�H�uμ����֔�����&�M������P�����J�G/��n��"�N�Ֆ?�g�y���a�$e˰�������ς$9�(^� F��cy��m���If��.�έ�p�l1Z�4+�f��B�6N�C6f$8[$���Qt�߃�X֯^���,DX���>�����vM,,�lr
�K�2�c�9�ή�ؽI-�Gr$����]����˰����?�^~�Mǡҙ����1%��b-��/b6@Y�'O.,���R��Aw�<�k+J��`�U�p�)�۶���H9*/�vݣ�u����ޜ��h����(e�c ��q�yA��3���j,͍��ko�MK7$Z��EBk�14�FB�:9W:�����ς�9���}��|@������B�/�3�������Y9��h���I�bcO?���^sa��f|o'Sj1FZ�x��7�m�V����x�*MMM8w��ªx�:k��FnN��0�<Q�#h��|Z�#w��(=�~�
�����j�e�[t��Ǟ���è��ĦM�:��7jpr2��SO=�pH>PKӁ������tOQ�w�}W���G�Brȗ��p��P��'��9rNc|X�ЍɅ��G�?��/�w1*l�eӌVA�~�m9�|��wK=ψ'9����u����(@N��Fӂs��j�<�b;�ӛ>_�|Y�DTDlj�ľC'0:�
cR��{�I��א\�m#��}Y�c�v���4��|����@�����_�p�����[{K�P��(��pj:���9�M+3�w_T)��g���r6t2��-�Y���-ݰw�"!݌~.v>�u&��oDK�Q�}�L��6o\����)�k�$:}��Tz#�׮]{e�6�I��zvk�z�]XBg!.TK�|ɒ%󺗅�����|Ff3&#:��s�6t���/�X���$8sJ)Ak�V�\>�η��w�Vw ++�		�ź�r�8��Ń"Ct-Ϟ=+Ņn��V)N;�)���)K�\�]�~��2_Ա��K�{��ъf�� OfT&%����?�{�ݘ��Z7n��Չ9�{���D�E��JEke;�ګ�T�1,���2��v�&����^�O~�y�^l߶ŋ�\��Ƃ�{�'���S�NIa!^����2�rm�2�IpZ�xcz�bI�|C�n�z����|hsG��7:G[������۷�@$t#�S֏�#��~衇B��(Y\���A\h?6�����(�!!��N�;����^�4LF�AN�k�*yM�v0��Y2n��/k֬�>��n���d����U#.���_H-�p��U�B��{;���r�CD�b	*؄�����Y��>#�R%� ?o��}\_��k֬nJ)"���߁������/�-��C�{��&[/�X�99X2���s">#���x���&2V����e�7�GG�[X���֎��c}��$��($4�Kr.\�Lg����,�(�|m���Eww::��;0����l�>��ɅP���m"�U�;z���
��2�U��`YY����|�H.�78	�����I^������+��~8�a����W�`L̑c*j���U��%��M�#����HN_�9���#G�eO�Pǂ~�^��t���o��.�6�����#�^4f�g�2r^3�)����R��F�����<rr�R�^3v�ݻd�%5%5$��z'''!3=	��U"PL/ɯA�Z�z�s�PZ�rU���
�����	�0���/�����}M�s��]��.[�T<�����wr�J-�������������<8�N
]�8�����'��Xd)�o~�w���Ж�*wC�������0o;���7��.���z߾}�����|E�y�O���+�_�ǯ���~��?� �s�2q���P��9��kH�'�&�hB׌��;�8����kk�74S�\�'�f~N�^xI��WL�[fN�c�.p�I?M��7K�۶l��������c@ljq�}���&�\���ƣ��6��}7n�%�p^��>*k1;��I($�
@�%֨�k�]��օ_3e&���BrӒ�����P*#xF�$z��Z<W���X��#����I�CaA~HY�i��=��#*���9�f)�ƈ�3�(?��V�Y����Ea�I}g.i3	�$.yO>��W�7������M����S�dgeN�X~o�\���R���<W�YEy9���C~�^�G�|��뒲�*�f�ox���e�
�����_jca4�!��� �����J0Tى��KH,_q�;:�9p���8X�gf����p������\��?CY�4�@S��g��Τ�LBEE%�iL��ڎ�v����g�	���_�|���<��+&|��~�O�p�����@L�&��CW�$g/u��`���[��{�r��x��oT��T���Ɠ�F��qo|�Wx��(���^�Ƣ+m?��~�����Ɉ�~�0�K�����k�W6�#w�,@L�&��C�)��t��c;�T1�coh����煏����0ߠ:s����/N�`��|M�~�7˺aϹ���l_���|0[�ƶ�%���>q����	�r�6�DE�<�<.�~ 6$���tYX�^ �p�'�Y�����`|On�;/-9���J����݂S��:�_¦;���>�~�l�z�7LMMFZb.��(h-f��2/�X�xg%o�HL^,��\Ř]��{�mEon��y�+W��C2�Њ��s���(dyV--�ts#��L&��N�l��IZQ���N���Z|1~����t �eq�U
|,y��6�tY�y�O;C�B�C�.��;��/B����O���k�����x���!����G{g�Vp���}��+��T2I<G�Y<�T �Y�UL*.�.Ӽ����2P��Be��`�
�7�_�������@�;H?�TL#>��zB����v�l��w�܍�K�cԍ(ux�froyC�FX�d���u":�&[��L%�yu`��.*��Ht.a�.�X�XcI�>�oGk�Ȟ���6��a'T�̟,�ght�������{���[(��C�$y(�W��nJT�p�OP1��F�L�Mܷ�f)6ܓ�7��PV���EAҟRt~G?����cq��������v��1�S&t������ZP�t]�v�F�t�M�a�j��M���A�j�m�x#�8��>j�4ܨ9I%,���k��<�L������O)@[�kxy�Q�`�8�w��d�����P���n,Y�|���\� ��G�����f4^l�,�3eLи��RLW��:c���EpB�s�N:tH�R��?!�i����I���G�}�I���,�/{�oo}i���<΋�۽0%�~$��N�3 ����d[�1��M��Dg0f�`�[��MmC���C%6�T���g�
��>�܃���Efx���E5	�(Z����������{b!r/Ų��'G�yw/���d�
�FL\u�1љ�Hθ`�g:Y��r��H&9E����#T����ɮ��)�8��) Z1Zڭ[�N��a@R�Fy���%�;�D��k1�AbJx�qTi��Kj��7�8�G醩��'�o>&F���8Hr�r|1z�ui�b�#�<����7rB��2��3��^�Ͻ�滰�0$�͸�޵`S�7������
�7ݶ;�3�R�|��gGG���
���ȴo�|tWx1�D�m!�_}�U|�ߘ��<��M@e�����[����%7Ԇx��:e�(��{���G?�}ּ��6���'�\�Q$$�Oi��s���}���O�sW���V�����b�ٟ�YHC7����>�{�-�m��v��MQ��L�z{P�Є;&<�A�6�U�"*{˩�I���؋sSU#q8Q~�ƒφ}���~)�QF޴�?��O�P3��&F�Zo.�G���c'Q�8����aN/!�@�� n���y^�شʡ��0���V�,�b�$�3&�
u��1<��SrG��/\���>,ٜ�~���~,���Ƽ9Iq��Q)0��� �~Z7�E���Xd1�'���	�j.����}^x���0���6֊(���,�P�o�f$�'�����hmm��%R����+�)E��8�amf�ڄ�-\N��K���_0���i�y�89�e�V}��c=/Q2U�?0���v�Uՠ�B��H(،�����bp�18p���+#_7�ݳE��ą��&J7��A
�d̜Q֘+��T�SOO/.7����R���s���W�'�نo�۲xp��i�IxZ<V	YD���Ҡ���h���bX�6 g�_�Ѷ��S՚S�Jé3er@;��7e�W2�ҍ�ϙZ�/�X�����\�����:A�E�"F=���3�I��������q���K_�R��I{��w�HƲEP��-�ḁR<(cmS���g*Μx[����E�-$�K/�$U��=&�9�>({t�b�y�X���²��M81)�i��K��v�]�����S	d���5s	*�Zc�Xi�2�c6�B�btkt��DP�(�I��{=@!�ݙ@�jZ��op:K��=̧i��1��/6nKG���F���\?��h�!�U�5�B��T���d���W^�֜l��?g*�n
�
�OG�����N�ӊg���=�5��8��jrԆƆz�F2!@�˸��t��2�j�S��`�9w=ʫ�PZ�II�!m%B0� �駟�A(O��7$83"tS(�ƻ�CY-��oF�`.X��cl��m'�{�!�]�Pym�P��ǈ]��5���P^f��aL��F6Ʌ%O,܈�7�Rm23��		��f`6��G��s��Y��	��D�gd2���>��T'f%7����9��;�t9�Ko�����܂�=�;�ᆣ�����\�^�T~����2��*6obj�?��32=��w��%���Y��&9�X��K�ĉ�J$&ąLr�'-!/zUU�lQ�~�TI3[ �Y�a����Q�n{«o����X
fv{��&���`�Aܲa5�޷QZ�X�X�+��c|����v껀����o��oe�/��/?�a�$'�b�H�[�֣ehlj�قP�6h�Itj��3�{�礏�$�l�Y/�z�JK�F�OGK�7��v/T��ǅ��5��/��U������S�z�#K�!T�EM�ߑ�%�7���ݻ�jժ+�v䓜D���6��=](+�ĝw��k�B�@�Dgj���[��"��PG��Z3fQ���e��f;��\ӹ	9��[�"W ��aJR���S�_���8ܹm-nٴq�ƃ�I�۬p�B��؄-�$zē|֜U�o��˫�n�j�L%[��7#���+��O�Ť%�m5\.�$5��ϒm$��u�&�l�hlj�Ɋ���5a�C�
q� ��ý�7���<��6lڸ�S�&�3��*�<'��)G�`H��Go=:���lYnټyʹo��/�~���?/�'I��i��[����X�;}��x�uY�{��d�<�i�nssN���1m��}-\B� l��H����>�իV���r�!��ƭ�^x�|���]8$'�2�c�7�?��/^,5��j� �r�ߔAs����w��O�mۦԱ9U����{���7��y���'�f�A녋58YՀ�-_�:L�$0�bﮃ��[�ן�P��3�&L��7�`flA��]t��R�}��߿�G����v��2�� �������x��7e��\b�q����=��f��?�f`Ř�V�Ӧ5��8xǫZa)�)�ۢ�4�f���;��G����$�p�m����������QX'��@�F�������$ass���z$�����KW���U�<pk@ta�B0�ś�~�dR��-��C�?�5a^�K0_�$7s�|���`:|�8��t®΄%kEX�im�5H�u����$�_l��;&��]P$'�<����Z��>�N� +����z�;�رcl�ޏRY�I�S�j�7��7Ƹ>��</�8x���s��<Hdf�:0�9S�yn��m���,z�S�J��
(��w������:b���u��,c��*�����D��&Xͱغeӧ>�r��e��A�2�N���'��t;�����!��R����q㠋C�n���\	��1�L�������F�SCN)��ݤw���b���ɝ��7�~�.� I>����V�����pY2e�y�� ��\���U:�$-<=Zq���}kZ�q!�qi�F__?N������(��?�����I�8J��M`<��]4�9`��[�
����x���ʊ�L��o{���֙d'���̶�o���N��3�Ⱦ��e+�l���0YTR-`6@����Mr),/.0�����ǫo���X��$�C7�7����3�P�b��!.�T�Ӌ�wۡS���;]p��j`���9�>��U{�]�O_�sԍ��Kd><@7�����8r�5.xb���N|�ٛ�a�<::j�w�[�$'�R�������^���s>���[�?��>$��cX[׈_{].#L�[��^:�%Fc��?v��ƻ�_A���\�Obωc������˴_�<��g~���2<���JZ���;�5%ݔ�B��<ΐ��>-�5�_`qˠљ��Y������{�ځ�+�����\��>8xH
<�
w���e��e��P��MB��-m��~L�^���:P�b�O�g���j�w�Uյ(]\�իVH�G��� VL�[Zp��)���gT�ٷ�5�<���l�]�(5gt��D��|Pp>6�*�}'��Ԋ��R.�� �
a����E�ֶv\�k@mC+�/�"�O�^���EsbKB�9�Q:tv�Je3�����g3���� ���dLƪ���@O�)���IdV���mC��"0M�R��m�����Ei���*Q~��(R��7i��Y�
���1!�����a;o\����d�Y!y�0Z�a\� �Kv��� ����!;ɀ-�7�֭���h��fˍ��b_{�:�s.A��+Fn�lL�Ot���x����v�6��/��x
ɧ��ӊoE|f)F{�p����1�'�.]��˗bIi�l��I���3�<WuU�ϣ��jS
`)D���B��W��,0����c��{���;�#9if�=<O�����SO)$�*�}�F�ZoG\�t�����e���V�ȉ2��jY���Ͳ��4$�o<XM�hX�)/�������������7����pjK�.��ޜ��uqirӹ�$	9�o�_�+�6mX7c�&<o��������e_PH$���I�N�3j�|�ݝ�=��[�s�H�
}.P�ߕG0�>�(�Ͱ��s���A4� V�8��
�(�U�0�4����ġG�����T�r{��>�A�o?FFŹwz1��bxT�؄��aḾޔ�h����SG�+��ۂw�������uk���˵d�������l��!�If���0J �'���� �0��@F��p�0jΐ��Zc��FJQs[qj&@«�FX�ÃJP�c츈��!�vv�7���%o[���z�c,�>�8�C���FK��xj�	1�hb)2��Z$?��J|�����d��q��֭FZZ�l��
oHn�����8 7��Q�$gPC�M%�_|Q��9�^i�s]��LߧR����EUM-2�݅��aL.�J��WC�	7"�|c_�-n��O�pl�������Z���󨹰��yN��7����	�n���z/ٳ�ɼ�믿.%�9o�mq����?A�q������js��g?����bK(}J\��$���9*���{ ���S���#6qf��H/2W ��Q�%�d'F�A<�t_��W�|I16
?�.'��U,�u��K�|�s��<��,}�kw��ؙen���7�)[̩�q�Љ0�7�]��c�jy	��@U�~xG�Ò�rN���L�|,�s"����O*l��a�A����	Cy�����uz�(1}mV���8}o�+�WHN��JL����"�8��e�G�tZqW#''[�;�8����aWk`H,���
\�L)0&��	"�޻���A����8?���t���!�i�i�������m�G�!����g(������oۆT1G��%�pL.M��9��ì`>a�m3'���j���oa��-��?��D[	�b.����c�=��R9ׂV�����|�o0�yQ1:���@�T�`^��MKQXEbS�?)y@=���!����������@�:k����>T�L��}�W���DwJ�;��#?��o_@e������sxd׭�ܚ��>�٘"�?�\��m%c�'S,L�Μ9#�A��	'B�R�M'p�l ��,l^�	|�/m8{�-��h�ۋ>�2���>��?����
��
f*��)bCg>��ޤ5ذ�A�ׯlB:���x�?�5^�<��K7^���X�n-��?��K��eZV�H��CZ�o}�[�M��r�����D�Ѝg���aPkҷ���(K�QQ
��*��P�����t������[��L��ܜ,�f4���N�,Ŭ�@��pBE	b�G}!�m���qԾi�.�F�qq`vl[��J&��Ʃq&=}6���� �PM���.)��X�&�5�̆K�՟����ay|=���X�I�N��wܻQ��pC5�A�ĕX+��,�1Կ���������h�߹i���7RP�TA�
�T31-]��,;p5�+P^�EX�	
Sl��#*F))�����E�������(���CŖEV=9�9����G�EEo��w�ޕ��F���]}�0XK����Y��� }H*�=gp��.���u��}�چ�ɻ��u;�Y����\1����;��u�J�P��@ņs��s��F$���Ƽ�ض��ZF��Ԅ��?����;v��m����47{���;06�Xr��Ν;���_�>@�Δ����#鶿���6�7�t��c��cY�t!*�5����A(�E�N:�4Hp����h�f"u�f(P0[P��_�~�����kI��������aXaL.��<
�d��sr�%�h?'�}��{��-��;��	�`JYe�Y�lB:ƴ�[�l�[�UTT�f��k��!�OS,����يsx�Ó��"!����%d�`��J��~r�Q��g�����B)��l�G��[x�����Sx��r�(gӓsB#[����R���?�~��`͚5x�ᇱaÆ�_�e{����gPv���U(��Ĭ��@���1�3o�=�U�?��?�رcx�g���OK+σ7µ[`SƂ�./����娫o�ۼ���`H�S����jv	J�U��$+����d�s�='E���r5���+��ͭƠˀ@�V����A���=�(�*&�Ȱ�e�ҥrj��͜ ����$z_?**�c$sr�I�r�}VLIyJE����eGf^X,�q��^�}EE%~�/����n���

�"�ں���Br��
"
�D<�+�x($W�PH� ⡐\A�C!����Br��
"
�D<�Mr�V��8#��{M����������Q�``Ǵ�ݜ6ɓ��p߽����,�&('��7c�Ӓ2�6�9��{���P�`.C��D<�+�x($W�PH� ⡐\A�C!����Br��
"
�D<�+�x($W�PH� ��� ˪,��{    IEND�B`�PK
     Y�#\
�  �  /   images/9eaf56c3-a2ed-4703-8e91-9b98c221ec28.png�PNG

   IHDR   d   l   ��9   gAMA  ���a   	pHYs  t  t�fx  &IDATx��}p\�yw{G�@�M�"H�U�Dٔdɖ;�3�d<Λ��3����$/��<�(�Grdʦ$�$eS;�
� �($Q�Bt,����}�?��� ��Y-x���s�����
>��`  ��A�%I���:���A$�#"�0]�5CRR����<k\�tww���]��X���Baz��g�ƚ~�?�B9�y���t���e��S �!L"���&�-��q��<o\�U�R���|!�L"�%��E����o��B�*|��!+k�aa�-[=��#f�R�jЍK	�L�1]"�l��b�JA���>�VfBc�����l��D�.�hA���t����V���6QT�(R9W�>��)w��}�__�GW[,�ߍ�(�u��͜���\�!\������h�����y<>�ٚ2�ɑ(v@��>-2���}:B�y�� ���v\�~W�\�>�R�Dr�O�%�޹�&�2���l� M��q��׆c�ZQg�A.�!�J`��!g/�T�.�f���/Fd�z)�z�h�y!�	0��3�w:��dg�߈��E$��M�;@�fT \���>7��.H�;�5�J	|N7Z{g�;��������ѣ0��ؼy3222 �� �].466��Qt�$z�V@�N�{FA+S�UbSn8�`7��z`Q����p�mv�4r��{���nD$�B��M�6���k�ҥaX)�ǖ��ӆ��fhS�؟�DS�	&ZډDH��a�2-�NT�W�v�ˠž�8;�����p`~D'HCC�9���l�_��b(�ref�/�kKY���'���)3e
{��csx`e/�ׯ�%"�K�P&���ϩ��eԕ6�D�Q)�	Z�
>=ՄzA���Ebe��$9*J[�i���� �F*H�z���^�r ';�-��J�*��/nEy������3��b���Ǒ��ǉ1輿�k�� �zh"�<��"En�8PRnF��)��HS�Z�nX�^N$�B���}���97��x����j�x`\�3n�	L��]nؙ�j�qs��rP��0�h�5m.�Y,�L$��7`�¹s�5�v������Y�lp��)ix����__�[�T�lq.F�R��%�l�l.~P"!.a�UL��6�:dgj��8$� ���o��k�(�#N�¥ZLj���)���
�{z!r����Nd�5fq�F��� 6I� �\9�JKK��+�@,�2��W|�_��~���ǅ�A�m\��=q	�;a�I�������@e���tHg��ɓ^�ks�����la۝�[cEk�%؜�ź4f�5�����#l2W���V��[���D�׌-�j,7yp��=�n�����1��>�����G�h��C)m6v��� ��I�����n��s�	�г9����ϕ*5��P~���TLdf�:l8|�������w徝s��i�ٲ>�h�A�Ɗl� zTm��j��|��lw��Y���,�27#깒��k�/9������$�Z��B��AK��3�/%��<��'V�LR���d���]�<�}�/KF�	��@��+���86�<���\�Â� ��G9��E�=�lI�r����.�*F������c�PrS����;��\��7n��ь�h����nŷaޗÐ��LQzD�]~a³��N��ގ�������G�t~���@��ޚ"��'�j�ؑ�8��q����J�����<x� 7n�?�]���+�دZ���(\_gO�-燦�F��vB�!��M�6������ͅ^�g�$X��7�l�Y2#v����/�<}O]���G>�c� ���<}�����o�>P4��ΜǡK��'o��T��n� �y��/���~���2�(fhgG;�?�Ck�&�T�����8H��.���~��"��_�җp��8p �W��*������Ǚ�
49#�M�
�R;�Ġ�Ġ�����a�0?V��/l/�'W���&tt�����I����S脸c�ҥ�p
E�o�.C��Rt�L��DoB�����C�KjN�g�O�]}���4��C�B,� U�ٿ\��ٸI�{<��h�����V$�d��1��ǟ��vjj*6l�����1$�رc��I]-��k�:j3��3�7D�@s�3�D����iGOk5,�!s�C#�C&vB�q0GU�S�6��[�@�>��^5$�x�cAe����af�8��v�设�$Y=v���W�N������gdo߾��Ě5kPXX�/��yX�)y+[~b̽5Er�ˮki�����=�H�T`��p�$�!��O��ݬ2�l@2QZ�b�Eww�����hv( �ʂ6&ru����&��a���W
4x����No:��K� --�W���J�o۶m��^��Sp= �����7%jĖeIX���;�:��[x�K���(��J��Z�EL�	Y�9��p�����(.+�݊r��@�R�bƸ���]s�����o���b��M&^{�5:tEEEX�uY��h�x|*K��L�������=�_D"йd�DE� ����rQY�'�^A��Rh�7CG)�I��9n�͖�$J�7�7!1 �&����.<��M�{��Ww�|غq/��9Ǹ=��"�_�YY̼O½{�q��5<���O̅�J=�I����.��� ưL������_X�+�Y%B�%|im6�[)���X��b". +W�d�ǧ�;�{��8ba�)�0�j��ZI/gf`� �N�%� 솺�A�zo�^���\N�,x�&&&������ƹ�/�������B��aA�F�(�������A�^&{��W�����>���D�R��w��,ˋ8v�s�� �OM|��#H�+>�2�� D����W��K+���.��'��Q#%�b�Ft��"�C�/zޟ��Q|�	�9�3§1��6�!������,^ۘ�%Kr�Iq?+Dyu�6�}xUw`L�,��c"n�)�h�������QVV6��	詽���2l`
��������F_��|y��s�$32"���X������(cp��]f,�����w^�
���>A��;_�ǻ��C8�dd,<�z��J�
:FD����U�x��9�V�>)sX�>�����+G��DzF��q��-�.�	|�obϺ��E�*e�Q_EEav�Hע����˃����q��
���3�gOX{F\�Є��
?�~�ݷg�p�?��j�޽���f�.����n�F�Ҍ��V��*�E755᭷��w����E��O��AUr��#Go0�pm.~y�.�Q��He+xF}\����;��_-�t�ld��j��ƍ�s�(s�hѢ�	��ֆ��jt����k�:��V��٣��q�\�/���LDDF�I�L���7o0'�˖-�]�RRR������/��2�ҁ�f�^~�2\�� �-�K���&� ����Pժ�_��A��8�M��!2*�F�K�����_�*G��Aq8�u�^��C�^6��
t��D�4hLK!W�݊@	%���z�.���i�TpA�{��yp1�ͅ��7��<|��YzK][�8� ;�*``��Ǭ�N��h�r\��-x�mлkQ�a���3��u"J A�!ǎ�X�b���Đ�r��ha=]T��;'���],uzD���jd����@`��	�t��e�~m��#\4��(`:�Ay�_l0�5`������V�n�Rm������,"����rt6���s
���w`�;� �>��!$ˆ��(�������[��~�Ƨ.�c3�L�Ѿ�GX�+�[VC�ycc#7������l����q���tuu!**j0R�>���C�΍��z(�atp
���y$r�)9%�$�B>��q%H���矟�����������ܩ��l�I&��8�c�L/ؐ�?��_tܻw����sY�B�".����I�}��h���d�xs���������U��B]�n��O�}��2?U���������՗V��@A�!�$C֌ F�A�1l����J}*ġ�?�
tm��,".��p���@~�<.�b�j&��7�/�gO�b!�:�q�W���&F�D꺝���{��綍����Q��}t��CH,��6����������![g�7(I�}����2!����ʣ
�m;�?�ي����f~򳿁�х{�es1��	G�Ѭ�Tܩ�.*y�t3A�s.p����ɀ �1�wtM�y�dm5�]��2�����*��:k��N����=��%֬��处8�����L䉬��U���ck�����UC,��]3�'C�-�����ul�v6�������1G�%K@�a���Z���炿�xb�t;���&=@���,�w�����EA����*t����l��C9n���F�fl�tu��#VL��`7���I���T�C�[���b��2�?*G�$��*H��/*�L�+���1>8p���O7�n�BX�:$��<z\��&��ŔT�x[=��Bd�5��6hԼD����A����|-,�@�w9�P��^y^���~�!~��"x�J�-߂o���o~ڄu�PEL�rLGȔ��A^x@~�%CAE�gQ2�cccG�+�Pfs7Dl$��g'�uh
�qK�T�����=V;��Q2�J!.�g.���p}�,��:�Js�%#�Y2T�J�n�j��:�ʝB>-̑��[�^��{ܳ	aժU�;%o��_�r����7��)*��ߜ)�.mה�C�&����O>䃾�����<�J!qJy�(�K�\[[ˈ��C���[�k��H1����?d���<���`�֭</0�7wu��ɳ��l_�R7�P<��d�X��� ,<"(DA>�(�J�s��uu��Y揥�z桎!��I�����y%�l�"܄�A���8�<>��#\#�A2��Q����\I9P%l����S�;3�K�ʇ5l�}L��D'������c��ğ��9��k����hokG]���/S/\�*lZr�^|�Ed$�QRR�,�n\�~��a�ɀ!i�&v�i��;��2q��l{�0H���$�$B\�p�/�h�Z���h��dsq5|�9�[��
D������D���ItPEtt4�5$PHU�O!��c\:|7гU���؊E�#���SR�;M�s�=��>��'�)73[\B�S\\��>;
�Gİ��b�����B�M�Sl�����܂�.<yR�x�#�GH���J�0c�G\�+���/���[HHL�s�.!QID9{�,�Szs&Ma�*��N1�iSځ��	B�����U-��n�Z�ߛ��jBWu1�>3LZ1������O�)���5
�0�������]�r\-?��u���T GAO"Y/��<��Y�߄�?�B�
��&���2��r1ZaB�1vJy�ۉ��D���]��_�͍�b�b�r�u��}ނ@���F��2 nmi�ЫIǥ�2^h@71t���ŋI��x3��7ȋ��#� �q��%>�K'B��{tnmM.��A����u/�p�Zw;�ex���#2*&�JߒYO��'O��ԩS<20���T.���������9KGx�4	�g�T/q
�jj�����8�d\��s�S]]�;�����HT��"^Gp�b1z��5�L!�N��bl[��w���8hA�������6o���t�E��'�_ßFF1}l�&��MY���U���C7��ǆD��v����a+��7YK��(����
*.)EI��YR���$/������׾7!1��5EL����wrc�������}�x�z�r��#� y�T�Hݫt��%
�RY������$q@D !�`׮]܊��h �R�����%m�R�����2|mW""��4��������)�PZy
��/a�����F%�
'�CQa�p�}UVV2B��e��HP!�O�1Z�U��ça3l�~���L[��9Y�����B���xU��_��r�Yl޴����V
�P
��WO�l �A
�Z��f��~g"C��'nlh���ΣE������9��w�DiE���Nw��K� ���R�����.����lz�a �>ÉEDD�����o-.bVW9����B�ɹ�2���C&�F�k�(L� B�EI�v\||	-���W�2�ċ�'*��=�C2Q/����S����}tZ�8U�� �P��n�p��K6I���zR�~��ؔ��5��3�Χ�Y+f0|S����7P�(�<e'4�hLw��@��ߴ;�h��E���#,� Vs,~{���}��kr��l	�#����E�d9"���Hp8�<Fw��M\��C�â�|��gz�@��J���S�"󜂜�����6�\V��'Zf�Ř�����g�v��f�"3#�Y[)P*U���U�?���"��y�<TQ���ʇ�({��*Y��S�8!f"NG�l]B�_>��["-}���W�1��{d�T��Վ>I�*�rkenR��H���#���BG[>+���;7`��G�)��0�*tZ���{{-����Ջچ4v��G�:	ڬ��������\ВwP���X�wu��������{�[Q���ݻ�	B��v��*�FI�J����Xr���)�J_�B5�;э���1vt1��rXلw�zG=J��s��a���⾈��e"H�\��/�r(3L�$�A*�խ�:��ջ�w?�%��/P�/^��������$���#+�B�� ��i�䮮N�T?ƥ��(*?G�h"�ݴ3-p��_�˂L� ]�_q��wn�����m���y�O���vE�?�K,��&%~��O�"�4�_�I	&��N��I���A�s'5�>|��!����CC�a^nBb�o؈M�%�������6&}63��9�FAjDLuSC&}^��⥵>�`7�p���޿{W#��mX��S|<�p���D�@���s�&�}<Pk�k��� ,2Ք�C�h�T�S�� g#�W���1�������?�X,�a.;�];���6~���<��P ���?���=k�?�����cg"������fJ ��s����GN�4k��
=��,�?�7�g��a�Z���5�SHTB�)O�a??$�P�Ⱦ���-{�wc�7��Q�9��b/'-��1嚄fq�p%���R�O��_�9&���_ݑ0��)���[��	ab��ޓ窌��ݯ�^���c��Ё�P��WH�N�P�!�Rd5�?f
�wHdI�I΀):�e	��Rtv�Q��Y,V�Ej=?d� P↜A�����,{.}�k������}��ه���/S�Hz~�L����vA�!
#v�O���?76�ůa��|Mٷ��������\�0s�މ�C�Fh@����((d���x��3��G �2yg5�S���kz'�Nv��e���#蒷��2�(\M��Su�/~�����`���g'�ɹJ�b61�2�j���!o���|���yK UtPe�T`�YPv�����v%���CM�����7����H[�����dɉ'x�����p�!�X!|²!�1f	#2�T\F/���,�����a|Ƙ��>|!15�7��Ke���y��7D���$�NB�\b����#D��	Z������,��?���0��0�1���S�.�=��	�R�Grt<��k�kr8�%��9�k��QRZ��l��&�i@�Î���|߭�0>ATj|�����b�03��玅	�:�E)B�����ABY`d�!D��� !modq    IEND�B`�PK
     Y�#\VX��<,  <,  /   images/5ccbe72c-6fd5-45d2-8118-bee80363f106.png�PNG

   IHDR  �  |   u:�,   gAMA  ���a   	pHYs  �  ��+   %tEXtdate:create 2024-06-16T02:31:32+00:00���   %tEXtdate:modify 2024-06-16T02:31:32+00:00g�JD  +|IDATx���ܗ����W%�0��
3����m&��9+9ݑt*�rH��N��
!c�&9�6�2��A�f(�"R��}Ws���������u]���Q������������w}���]I�$%ʀ%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR�X�$I	3`)��I�j�Ky�;��f>G��a�R�-�ߌ�C��H�Tt,��8~M3�Ћa!d�A���2`)f����6WЇ۹�g�$�hXʎ:�`&KV��q��B�s"Q�^�.I*��c)oҏ���E��ڭ�����?
m��$IJ�KY�Е3��,��W>�>��Z���Rn�j^E����-K)�n�BF�?������F���$�.��NB�����=�r�чn������ ��J������&�)�$U�KY�c��p!=�U��o1��}5�|������C��j1`)��8S�]9#D���`�jV�͹�_���<�$IUf�R}�.µ9���ϥ<��kܶ!��65��;]\G�T5,e�+������1/z��B��Pn�#$I*�KY��J���4���r�0|%�M���0`)��e�Md��9����r�@��H,e�.f|b����=�nsIR���7�N,Zu�3n�4� I�j��EKY�άϏw3.�na(� I�*��M��Gsq�Y�!������$IZ	���C�aP�Xg�b���80�ٌ�|�$I_c�R���>�����J|�f�&�=1�8�}�$}�K��iAiCW�H|�oH�М�]��,�ŔКQZ��Ǯ��}6��\$I2`)Wfӛ~GZ%>v3�kna�CI�Ky3�Q��-�hG���^���CI�=��h	�Bۅδ�Q�W_b�CI�/���:q's6�I|����o$I�c�R���@s8�b��Ƕ`(I�e���M�КnW�wĊ��(�G��,i�it���2�CE��B&X0���0`I_xy�4��!���v:3ʂ�$e�K��bN�P��C�`(I�g���i�4-���E��aE����$e�KZ��t�rN�[$>�CI�4��:�q�e�Y��`(IYc���d�4?�[Z��9���L$Ia���<��q'>v���f2C���H�Rπ%�{������{��]���� IR����,b\hm��Ex�4_~��^@��Z,�*��VQ0��F��]q��i%)�XRU�`8��-JR���(n�p��;o�`(Iic������&%)}XR2*
�8�s�9�WGp=!I*y,)9��`8�K�����$�����U���Y0���2`I��2��[�� I*A,�X,JRn���(6����0�-JR�2`I�7{y��<�����
�3i�P�J�K�_��^⣷�,�~IR�3`I5��ît�`(I���%մ������%)�XRm��Q��`x	c�+H�j�K�=��8�(��-JR�1`I���î����
�ӹƂ�$�,�T��[0li�P�j�K*+
�e4M|�e��)�a��T|,��T�q\�
���VQ0�B$IEd��J�|F�te%)�XR)Zʤ�,JRJ��ҵ�`؍{Y��E��`(I�3`I����V��W�*�����ҷ�`ؒ.�D��G�(v���1$I�0`Ii1����Hõ�ehNI*I	1`IiRQ0C���Q'��W�a8���$U�KJ�%���F'6H|t�0����t����������0���\�H�
f��ҫ�����L���$Ā%�۲����Z��ac�8��!����H�"��,�Io���"_bths�$E0`IY1��������a<�$iXR��(v��K|��(m*���b$I�d���g&ݸ�c�A�"��_ho2�a�A��R,)��[0�}�����g�$}�Kʮe��ũ����h�4�2�ϐ$}�KʺE-�f,��E���Kʃ��]Y0����I,)?�]0<*4��Tɀ%�˲�����m�0zE�p72�7��3`I�3�r��`�)���݌b��S,)��(cJҵ�G1�����1`Iy���b�aXQ0��˸����$�Kʻw�q$�}zq�Sn�PR��$�(6���&>z]�i��&"I9`����,zs9�s6�-��r��`^A�2΀%��>bThm��E���~���},E�2ˀ%雦�֌2Nc��Ǯ����`$ׇ8'I�d���r��M_���W��[0�K�5����9,I��	�BkM7�+�O�&���,J� ��5�Fzщ�|+�g1�Q��$e�KR��З����S�ћ3���P��$e�KR�EL��`x,��1e�M��;�IJ5���T{r]آ���lF1��HRj�$�m2��)��"�ތ�e"W�/$)�X������2��(���Q�W�b1��2,I�1�N\��tf�"�^Q0|���=$)EX���r�ҵ(���Co��j��$��KR>���v�Nd��Go�Q�Mc(�I*y,I��'��IG��MFo�X�_�xI*i,I������ҍv�I|���E��1I*Y,I�[¤�ZҙSY7���^^0�x>F�J�KR�L�q,=hU��[s�r##xI*1,I�4�Q�)Z�pSzq.P�$$���$۲����JM����O��&"I%��%�f̤7�8���T��w�:2��yI�u,I5g~�2�QƑ�K|�Bx�����0K��Zd��T��V����6L|�����\� I�Ā%�6�Do�r4�sFo�.al��e$��$ՖOZ�rD~�_Y0��P�`(���$ծ)�mNg�q�c����fr=���TcX�j�[��?�Ѓ]�0���B&P��HR�0`I*�*���Ʊ�O|�Ɣq:3�;�I*2��R2���$��;��]��`��C��$�KR�y���p��oFߎ��[�sHR�����6��9�Qh��`��/b!�û�Ɍ��B|���ZSF&>�za�2�R�],&o��2쳛��6f,��¿�����Ϋ,AR�����6�s8HU��pȚ��<��sxH��it�b:r[a��B{���"��bO���_[��7Ƣ�=v:��o#�@,���A��:�ݩS����v`��&15D��К�wy��,��'os�Л��ϐEu�!�ȃ���έ�j��B[fv����sD����8�О#��n�GZ�2��\�f4fEXV0ܝN��:��� ����P&d�ը�!�_�4M`�f�%�%!���񼆤52`Ik҄����A��Z�9&��Cp��fO��Ջ����E�5c�(F�.i�S�c;�i£�e��.�/��V�*�Vπ%�N:�xը��д�������5��r�ю�E����U�ap�~؛:�c�n�kC���LE�*��UiC/���ڑA\���r�K�7��!��ʺ��ހ�B��8>!M6�K�I�׬Ǉ6����(��K��:!X]�^5������T�Q�M�f��Vy�a7�-�譹�K���Alʙ��I?�~����&�t��΀%}ݡ�S�wk��!��Q�qi�(Vۆ�ծ�M�B�����D)�0D��"�Iޮ��\��H���e[������u=o�%ʒ�)��T:<���]Y0|�����1��'1�o��ؙ�#��t��j�KZa-��2S
6e,����\�ͤ7Wp,݊r���!`]��,�)
Z2��(��P����H%��?װ�d�b}Y���cchKGR/��7��q?�%R0\�KB�,�����'�˟齅R�RzsJ��=�W�Cru���r4ϢX�
��qzh&>z]�E�et-�V��Δ��y�+��ϑr΀%m�x~D�jœ�O9*�K��r���ܮЊ!\�X�
��#�0AE2�ҋ=9�� �Kyw 7G.~[[��yk�d*�G�
�]9�?���va2Ck|�F�1O���3���B�KyV�K�0����}�X��T�)�mK�I6J|캕�J�`$ׇ8W3v�ZQ�����K�V�e�R~��u�BZ��T~���U�2���1����0z�� qk���x/�ccҡ}i�a�Y>[*�Ky�9�4iʟ8�?��Xĸ�ZӍ��s�	e�V��a���49��8��H9d�R>5�^�#m��n�`��it���\��9�g��g�\O}��`&ю��rǀ�<ڒ?�Cb������r�Ӝʛ�?�a8�n�f�m��v"�U/��r%���З����S�ћ3���P��踽�sNj1�Oy���ٷ�;�%�{lE��(�fa�mI��J�{���:R���?�?�<��p ��#LY��Y_��Z|�i���o��6U�"&�VQ0<�g�S�Tʹ3�����F���+���8����_���X�`�cx������f}�f�ZR�y�w
�f1O�68��ZsǱY��A�ˍ��*
�=9�.lQ���mv���s�9ҩ�����n�o!q�=�
�b٦�О���ݶۆw�!�I9b�R�4�v���/0������b��'?
���W�e������>T}o30��)��"�ތ�e"W�*��3���9��CH�C�8�V�odKNq��D���CP�)7Xʓz!���[�9,��Gl1���-΢Ti���=��)(	�./����(���Q�W�*�}��L�����m�g�)ͽN����*_����/��/ ��Kyrm�_5��ǣ$�]�2���Z�5�q7��<J�4:q'ә��0zE��-F3��;��U��aNt����b�Ƕ\~U��ƙH9a�R~t��#/�� �1�K�Ϊ�R���՚y(9�0��84��b7������kT����Jg8�p3=�}�תL�-#�T.<#�X�QN��;�g�>f�|��t�FF�w�[6g4Ǡd}ν��ʙ�X�i=pTh�ʄ5�q~--��O��OR\��%D��U��p��i�0`)sG��y��̦&�������XG3)�,%�i:�3���٦��flx�ǆ���*���	��1�qK(�O���]��-p��!X�Qc+7J�Ȁ�|I��X~���:jK�ml_�vC��g��C��^Жn�Kl��/lF/zpwx���0�3W<������� ~�EN�Њ1��y,���X��ѡh�]��?i�uW�6�=l�joŲ�����ũ����k//�b<����j�g\�aM�4���L�&6-h�cx��2΀��ۊ�n�?��\W�1�����ʂΗlO?��b�A7.�X�'���*b�e����-(3��KȗpC���3|ٱ�m�C�z)�Xʾ��<<I��݁�7���,��9��'*�y����`�	�87��XZө�mS����m�'���n��S�)S��0`)�~����T.�\�n�.G���u�]#�6�ݲ�asN��i������Mڱ��j���U����!x�;2��R���m�YP��8�$�~���E�߃S����̢7WpgUi�5٭�����Y��ka� sK�z���^��9�0���|��{r8h�B���W�~D���yՔy�]9�
��&�3~Y��bN�	?����)�Xʲ��Y@ￇH���1�S}��\^��;��)�5��ӫ��Qu-��t|�Q<B������He�R�]P���+��oa�fC:����j���r4�s?rwn����P��<�wC��T�(��k�f��$ K��6�]�ٷ>=�j�'���`xD��T��a��w¿���Ku�r�kPV��]=Y;�o�����#z�S跚�WTl��)�,6.�cU��U���;�"���W���I,eզ����Z�Eh�pt���pu�Moї�Cv-�T�q-���G�?�#�vb �A� ���W�K���tJ�s�{�6�o�ppծE���t�؂&��׭dϸ.s��]Tφt�|�2`)��pft��%wq�׍�=�E�\���J�4:Г��+�G�R�s����Ⱦ�Ç�yH�c�R6=�mL��-���<ґK�ӽd��@s8�"r��t	{D��#��\�I�W�%z��Xʦ�+@�䚥�yQ�V��GQ��������4L`��/�НG�E�ހ�,2`)��!#�e����b�eӨ�X%h��kؑ�زZ��'5���A?�G�< �c_E����=u���W�J��iW30��/�R��Uke�^���9e\�1�*��n��[��rW e�KYtBd�߰���yQ�+5�p&���Ye�p7�����8�0'z��R��r.��y�K�c�R��I��~���U��oT�X%�t�W�=غ���K��ׯ>�ѯ��H�b�R��ox�n�9QwG��!����A�K�hGW�,i�+��qV���.�0��,e�K��6�גT[�y�[�&Em�><�J���c�]tB(K�k�M��~r)R���5�gT�ɼN����u�@V�4��7��y�Ǣ>��C#>F���f?D�K���b��4��w J��s�/�g�h|��׀}y)CXʚ�h��;I�������b��]�_����~cS0��LdXԄ���-,eM�ـ�R?n�
X�i��j���� �F:-�����ΕRÀ�li@�~����o�yD�}X)�oT�7x��z8*`}���)3Xʖ�"��ɤ�#Q��D�7k[�oZ�{��i��)}�K�+^�%�ˀ�-q�T���`��~-X���%�`���W�ϾuY�J]]����U���G��C�2e�k@J�G��;i�2s�h�����R�5#z��+��ߣ�!aߖ��1�Y�V����H�4�t�uatKV
ĝ�I��@�oS
����%B���-.`��!T�XRF��?R�HΗ�ĘˊU۶�����:Y)WXʟ�)��q��5_��ڷaT���s]�,���+,�ϛ�]�w`�J���z�Aڽe�R���?sI�9Q���ҷAT����!�K��>i�AT����U�D��{�KY���@,��"�^k���*��M�w Ȁ������[7�܈jW\�J�"�,�KJ�:Q�\('��h�{�KY]��1`)�_:�;7�9�4�;7�v�ϻz>U�c�R����FQ��_Vʃ�܈�[�>+e�K�7�c)���j!*}G��(����]'Ȁ����ڱ����ϝ�q�R�'�M��N*�K��5i�MT�wQ�;3�5&ݶA���g[�N��I-�z������Z�n2�F*�K����iw���J��Q��"u�jN=��1`)�Z�<`���5���W)�/]i�R�:`M���vʟ��+��z4��7�����"�ꟓ^qk]�2�3Xʖ���~���Q3y��5X��.s#�0X�]x��j��s����%�G�a�_LZ�����������ڦ8`�e�R��-q?�Ӛ'I��zy�J��Q�@�"���IT?�Ye�K��:�~��ڀU?�l��Q:<�k��ʧu=¸��x)CXʖ%<A��~�0�tjúQ�G��J5f_#�~��q�"e�KY�hT����
itbT�I�%��2�� ��	)X[G�s���),eM܏�:Gҧ!����h�o�ϗ�y��F�;�n�KC������L1`)k�fN�ҸS��`��~��䑨��$����;�:�!e�KY���CY����H�����t�}�:�0`�9���+e�K�39*`Aw�']v���~�Fޙ���,�qD�����"��#��	�9,e�]�ZZ�h��l:��#�f���c���ᔈ~u�MGҤ9GE�[½Hc�R����Q3�ԣ'���8.��x�.��%�Lz\�Q�����Hc�R���ڰ��*i�;���*SP�<bӶ��s�I�����~$P��Ew0<jA��\���K+N��9�a�,�.��y
CRS����Q�p'R���E��}�g��ȣ���ȃ܌�g,P'�_��'��4h�	�=��#��1`)��G�:g���vm#{��%sSi&gϨ�s)uk� +X T&��M��E�܉����ք���^����Ȁ�y�����|/��,�hP6��M�3�Q�}���]h0�G�|�aj��ĭ�z~'|$(�����X]�I�d�RV�ȯ#W�1��XH�:6��
�RP���}ƕ��{:��@V�2�u#���8�L2`)�>�j�D��.��Di�>�L�b��k�G������y���w�"e�K�5��$�o��Oݥ���qt�+���'�#��Ⱦ��u��E�i_�׷�)�Xʮ��puEt��y�'(-�����{�)�\�J�HzF�JXaWn�,�������j?(�Xʲatf�Ⱦ��;Ji��:\ˑ���لRo���g�(�����]�0��k!PJ�e�R�}į�=�wS��~�B�������`�	�9�]�{��6}([�6(��(��2`)�&�����ޛ���Ȳ��"�NYf	�J�X��XL����.#��l�ClY@���)�Xʺ.<[@ѢOr��v�a =�����a*7rr��=BĮ];�`A�jQx�R���u�����
��m�� W{���ê0��Qv����K�+teð���h{q_A���f�j��Xʾ�G��7�O��NjǆL�GnӋwQv���=��8���G1�Fm1��Hg�R�}���:�.າ�����m�����-�9��;H�'<��?S�0(�S
�(<�R��KJ�Ky�zE��B��h^���	�A�]�V���Piq*����1�qi�^��u�@�W�[��SH�g�R>� �(p��C0;�����#8��q����cy����}؃�jh����>4)x�;.�K���Sص�����:�7��~x�~���~�y!*���������{����[�I�Ta�W)�U?����U9#P�5��2�bi�`��Җw2e�`�goՈ>G7�X6���Ua�E���H�`�R~������oW�.�����ğ��\^�kX��{�~�eKCP�T��D-x����;��ڄ���Ba��:x�U�a�R��ʦ_�̺t��1fvBϥ>Gr߫���9Ե3o!?gJ�o���<C�Ll�����0m��u+`�*)�Xʗ���:)gC��6���T͂�N��cx&U���ʾw8��͑�e���31�S�u.k}��A,��M�1)GXʛC�)l���j� ��~��m��� u����I	-J��z��x��E���)e��b��<Y���[ӖC�3��y�eƔТ�R�0`)o�҉�y��h�ѡU,�3�'¡k�Wӻ.[ђ�Áj��^�^�%�&�+���W�.�/��š-dj�g�
{�k��~�q�cw`���nG��į�J�K�������$.oZY��d:��.s�`����Y8P�����/�C;�D��8s_؟�k~Z�O�;�����/�j��1ۄ}�;$��.�)gXʣŜ�P�%��$|HZ��k��E��W��A�Jl���ZMJw�^)�Xʧ��e.��0iCmz>ī�Q>���!bU���ڰ��\��K,��P�p�I�'9�;s�?��І����L@�)���ffrې�9��(����+i��2)�Xʷ��7Ҏ�6�N�	P�O��c\_�ij�}t,��RR
��w��S�re	�
��f!�p'�r;�R�ӏKW;��,i)���[�C+9K��O����>\͙��W9��"�K�0�9��Y�R2�.<��M�Й�B�މR���\�<$���З;��a?J�B���箴��[�Y���aJx6��&-g����/��d�qm?���;���3��}�uxm?ޡ'�PT��K����6�zq&�k�9��K�R�W�9�Ї�k��g�xI_b���nnX�B��Ɇ5��SȽH�y0�6a�=��yׄp5I_c��Vf^:#85���k�1'q1A��)������N=⻌d���7��,iU>�������-�o1�y�z��Oٙ�Ƿ��8�3�����HZ��:���I�V��?��p�z��H�x�s8�}���r��L^A�j��5{���v��	�k�f2�.�#%mIe��<���a��,�1�7��FR���`]����v�b�p>O2)����]E6���A��=�-Uq�ٕ{�C^m%%fA����-i~�
�կd��+�^`�k����fThu��ڪr���}�a볰�a���<�RU���y����Zl�&ᐵ�h~-�:̩lo�_Rm[�ҋ����ؼr��ZM+�f!���r�}�׽*P�.�T}�y94)=����2`I�$%̀%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR�X�$I	3`I�$%̀%I��0�$IR���'O-�@�    IEND�B`�PK
     Y�#\��s��  �  /   images/e4bf1f14-66df-463a-8792-8567b691137d.png�PNG

   IHDR   d      ���   gAMA  ���a   	pHYs  �  ��+   %tEXtdate:create 2024-06-16T02:31:32+00:00���   %tEXtdate:modify 2024-06-16T02:31:32+00:00g�JD  �IDATx��kHTQ�?�)�OP�#��
�Q��BȂ""����B��V���0����bR�z@�!�C�dDjTD�� R��f2q�j�{Fb��^�{�e���^{߱� J$�%i0!�D�q�OD L�t����S�ijd��#�#����9�-�4��Fm����s���
��p�����~����p�V;��f�I�Y�3N��f ^���W�IR)�D��WG�*�H�4�J�*�N��bUj�qHѮ�(p�~E8�g:c/i�o ��,c�8@���À������:s�6'�`�2�-�*A��{�MJ�%y^�:�J*�E`(;��h��&�]���D���~��F>qȜ�$P��fd�D��8�Y��,W��S�"�w�bFd�h�Hp=�^�zNv��	_�S�I����z���lߓj���}���2̈��,�<=�l����e�/��#s����$�mFDb��8���a,PI���Sy�ϕ�:\�\�ssS1�+��	����]欖Pz6��>Z#���=�7Z��6������fay���1	�s��^�������i�yĚ-mv�V�¥�7Yu�o�K�nˠ`hҬT�����dmA���e�{+)W����,��v�ѧ��f�J�*�*3�y�����[��%��S�%�q�/VV��o.n�3�����5"cT-�&�w�g�ʐ	��`�}fHf��/T�UX��^0/Q<:\�V�U%&D��4D�D~��I�
��    IEND�B`�PK
     Y�#\q���W W /   images/7c9bed20-c7d7-43dc-b689-820375f46db8.png�PNG

   IHDR  �  r   5)�   sBIT|d�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<    IDATx���{t��}������u�,K�,Y�K�6$�@�!�����4�%cH3�c�$�==s�G͜�4�9I�`;&�!mN��j�in��K�IHq�p3$˺��E�m����?d l,�'m�_k�%Y���1kyi���o�    �wy{�����B}.Kf��L���Um��To�jIU���^c��K3%%�L^#I.���0����r)/i���4��_�#2;t��O�u�h�ȥ���z0HC.�4���>�A��!�=��ߓl0;�9�,r��4�C2X[�����7��      ����+WU���+<_��bMII�BZ
fYM�P�e5&+X�5�� }���5~�ג̽���_��L��ߺ����rU���ܯ��
�^��_�:�[kX���ˍ>�Ҡ�!��d�2)5�I����on�|@���>I�if}I!�5����u,y�?X    ��b    e���\SSScP֤��(͒7e!4ɽ٤F���U/�,I��jcgOaC&fR�������i���������2;�I�-�,)�4wp$9�I������c��       �ޚ�V��$��4����nu.�s�!�2�u�LIu�>��je�)�L�kM�s�BG9��l@������}A��-y�{�ue=�vg
=-���(   [�  ���zݺƴ427UrJ4���� �u�)��Hj�݉�l��r����t��{�Bo��zf{<xo"ﵢw���ӱ�?v8      ��a^�����$�l��l�3�F3�-�F7�m�f�T+�L�f��I
��q�L�s�S��2uJ�ky�4�v��/Yf�z:n��c�   Sw   ��_S�/j~b�*��2͗Fo.�)NZ����}�>w�YP��vɽ�G���\}!�]�������Ñ�      �ym_�*f�s���T�z�T/��nj�L�f�����FN��4"�N�v��9���vȴC�vt�����۳ؑ   �d��   �N��k꫊vFf~�Kg���v�LgH����AIݒ:M�+��i��$Sg��d��ù���߸�@�P      �ܴ^���X��ZB��$���<�7K�d�l�ܚ}t�L�!�����&{:�=-Ϟ��t�7Wtǎ   &w   ���mkOJB�P���A�u�FOao���I;%�-�r�2e/ʭ+�l��v�;w}{�@�P       ��n��r�P�\�\�����[�B����u��I'I���
�}.=c�S�-X�M�=��q��y�8   `�1p  ��Ww������+���,;W��&-�dL3\zI�n�~-��z!1��S�U���Eݵ�;      x��6$IOk��TSx�����N�L'K:I�I�cg�ߥ'��qW�.��L���X�;v   p"�  `J��~M}����ȃ-�k��s�϶��2�OҎ#7��w�n���C�������     �i���5����[�|�曍���*�4I�q��Ϥ>���|�����oݽq�vN{  �T�   �V�u�GJ�E��"�](��}�X c/��)��_pٯ��7�*��М�ya[�ґȍ      ���6$��:�,���N5�i��ͤS]:U�<I�ȕ@Y:<zT����$���{:V��   8�   �.oϵ�n<�C�ăs2;0)uJ�&�w�iGRʶ�����~�^�     ���7��id�/��|�1_N`&�Nwm5�&ۜ&?������    �B   ��ᣫf&���`饞�e2] �2v���(�yw=mf�����?J�3���}Q��Y�@      ���ew�*M�H��p�3�~��ΐ��X/0U�$���2e�,}hw��=��   0�0p  ��hi[Ք)���/3�e��SR�����Y����s�BxƇ���+�c�     ���]���"�s<ՙ2;#Hg��t�ΐ4#v�q璞��!s{����{��;cG  ��1p  ��h��Wk�ʡ�%-q�ȴ@��	���H�M���-H�=���}�'�b�     L'uׯ�/}a�-��B�-��@Rk�6 ��i���ɥM�$ܿ�影�   P~  `l�mH��.3-1i���$bg���������k[�oWjۺ6�x^2�     0U���g��o��ۂ̵Ђ��6� �V�vH���&��������I   ����
  ���a��s�}ȥ��~� ��^���|��m�m�R��ӱrw�0     ��d^�W����������/�47v��6$�-�/����q�S��   051p  ��;|J{0��d���gJ ���ɷ�m[&�^SS��_�q(v     �xk\vGk��E.-r�E�Od�� $=/���;������o�  ���1   �P�GW�̗�t�Ur�+I�c7�1��]�c&L�+����;     �h��WkC��yJ�;�]��N�ΓT� �A��Mf��e��������A   ���  ොt������g�f�ߕT�	 �H��m&���[w�����۳�a      /=�=Y ��l�\�$�-)�n�1�I��K�V���x�3��   0�0p  �$�a�ꓓ,\-���t��$v L��r=������,�Gzf�'t��b�0     P�����'��J�p��_ �&�SRC�4 � n�[3���4�枍�;   �1p  �ƚ�V��Z7[&�"��! �lH��dz��	!<ҕ�~RK��a     `�rk�f��!I/ti��.t�I��� `�pm3�=r��]�\�   ���	  `����/�*T>왵���%�b7�1b��oq��P���}R��Y�0     0�4.��5��"���"3],�1v L!�]�[��{�߶+v   &w  �i��<4���p��_RE�& (\�j�G�푐�#]o�;
     L��mkOʅ���Å&]��cv ����#�}�S�b  `|1p  (c�׮���o��ZI�b� �4�W�Gd��+�I�Xz��o޺'v     ��jmR1�;R����Ã���� `���[��k���l�6  �w  �2Ӹ��$m.��2�#v @��i�f�oɤ�s���mKGbG    �7�|͚�����Z�E��-)� �]&�{y������  ����  �,l�P��h�n���$%��  o�d[M�c�~��?��X�;v     �]��k��.6��$�X�E��1`*�b�w�r`}����P�   ��   S�춵'�?��Ҥ�c�  NH����FOz���~䅯�8;
    ��ն!iɺ��r�H�K�Z,�lI!v �-; �z)�����b�   �a�  0մmH��烒-w�J�d ��a�&�G�m�����+�cG    0U5|t�̤��D��ʵ�LJ�� 0N\)غ�����o��  �c��  `�h�z���&�>)��= �(�2���l�+��{�O�    `�jX���|��>z:��2�+��W��-K�vu��|�   �9�   �\cۚ��[\�IIU�{  �J��~*�f�o��O����     �U�5k�{�ktоX҂�M �I%s����wm�eS�   �>�   �Q{{h�>������!�s ��HzԤ͒o�{Ŗ���;
    �1wӺ|c_��D�Xf���I��  S��Q��TUS��/|�ơ�9   x5�R   �HS��
v�I��uF� ���Jz���<<$���X�;v     �k�G�8��P��e�I~�d�$bw ��N��$I�]�,�  �Q�  &����sv1o�Iv��ٱ{  e̴C�˴YJ��q��     x���UMn�Œ]"i�K�K
��  ekX���e�gwu,�u�  �鎁;  @Ds��r�ґ��{Iu�{  �R�I���dY�e�ƕ�%��Q    �饩mu��]�Kv�K�� �(�������q���1   �   D�|͚�J�߹�&I��{  x��&=$�-�lsoǊ�1x    ���ew��'���D�Œ��_ &w�wC�g���'�c   �    �@�׮=W���5��t SC�\��f�@�9�W{{;
    0�4^{癉��\v�K�3���M  �M���=+7�  �.�  L��׮>'���\�KJb�  pJzإM��Ի��Q�    ��z�	�ҿ����M  ��-!���{���  (w�  �Q�5k�{N&��Ű P�z���L�ݵ��c��$��Q    ����A���$��	 �q�%s��ގ[�  P��  ���k�<3���d�İ 0�x����d��e��ގ[��]    {�V��s�_
���b� �fL�nB{�����  Pn�  �����5�i����)I��=  ��]&{P�[R�fNx   ����mu��]z���Œ�n `2p�w��O�l����-   傁;  �h�誙I1�'6:l��� ��e;%�ߥ�����]����E    ���Ҷ�)���u��+$��	 �I�(ٗ��>�}�'�b�   Lu�  N�M���}�n�ɚc�  0�vH�$��4���c�K��    `:j���k4\�IK$-q�|I!r  S�!�����u,�;  `�b�  �5��Y����\�c�  P&\���t��_̧����bG   @9�����bRxo��+l��%�bw P&�e���]=w���1   Sw  ��Դl��������-  ��Ԥ���އ*��?;
    ���I�z�e�%6zJ�bI���  (sO�§{6����!   S	w  �ct��w�.��/\�RR� �i�d�c�6I���n�X:;
    &��k��W�������f�n `�ڔ���y��'c�   L�  ��M���}�[��/%���  G��c�6�kS���G�ޞŎ   �X^3h����M  �����������Ď  ���  ���k�\i���tf�  ��H����OK���l\���A    0���>9��
3}@�+$��	  ��N�������u�<v  �d��  �(�h�ܐO?'��b�  ��ʻL��\���]�=�    NDK۪�4�.�%�ĥE��  �[�z(dي�o�;  `�a�  �J��yۜO���f��  cȴC�˴��������w�N   �7�����h��=��HZ����B�,  0v�&_���CO����1   �w  ��Z�־;�I��c�  �q璶��~��?<\|`߷>�/v   ����uեJ��Bz�g�~�I���  ��yW��g��ߋ  00p  �^}ۺ��e�Y���G  LW��?���٥V�qb   ��v���*�׆�Lv�ܮ��"I��]   ��YHo�]ۮ�!   11p  �Zӵk��k�I'�n  �Jj��%m��)�C[vv|z0v   �)�mCҨ�w�i�\��t�����  ����\�ձ�˒y�  �� �ii�G�8�PQ�9�n��  ���I�����`�g��p�(    �_�5k�+h�LK$-q�>v  �
�A���=+��]  0�� �i�y��\�V�I�[  ��5 �G.m������úky1v   ��^9hw�
I�c7 �)k����,����۳�1   ��;  �6��^;�����X�  Pv�%�ĥM��Ի��Q�p   ���ew��'����]W�tr�&  Pv�d���v��T�  ����  Ls��^-�$5�n  �B���i��6�v���d;
   ��kj[ݢ`���D�ߕ���M  `Z4�?��e�5 �r��  ����6T�7�n��  ���&=$�&)�AW�m��   plZ�V5�!wyp_,�%.] �g  ���W��7���mW�  ���/  �l5_��bw}]��[   ^�Ӥ�rm*&����W�;   �����3��Œ�HZ   LB�r���c�7c�   ��  ��u��}i�I&)��  �f\zҤL�`Z�����坱�   ��b^�W�a������z�L�bw  �����P�������  0�� ���x�g&�ΥE�[   N�Ӓ= �i���X�R�    �\�^���T�.5�.w��$�'�  `�2�0ˮ�Z�ñS   �
w  P6�,]{��_�4+v  ��4i�\���]�=;   �*Z�V5�%Kv��%.�/�  ���$�l���Ϩ�=�  p�� �)�����n��  0A��-˶��x��A   �d�|��9�g�b�~�x^  L�������Ov�  8<�  ���׮>'u� ���-   ј~%�.{�ݷ�v��T�$   `�4,[}r��e��R�]f�9��   ⱝ��u=+7�.  x�� �)kε�����H���  0�t��2m���9j�鶎�#��   ���|͚���Œ]"�bIb7  L2%�?۽��3jo�b�   /�  `�9톻+׸tc�  �)⠤��9S�`����ΎOƎ   ������E��K$�L�Hj��  0E�c���񉽱C   �w  0�4�Ѫy�\n��w�n  ��J&=&���lsa$���o޺'v   �zպ�be�����f�TR]�.  �)��Y�������!   Ǌ�;  �2���^���%5�n  (3�\O����m.����w���Q   (-m��\����er[,���   �̀�n�w�7b�   �  `Jhn[s���On  L�Nwm�i�ܷ��T?���n�  �)�mCҒu���l�4zB��s�s�   �tWw]r��Z^��  �Fx�  LjMm�g�W]�4v  �4W4��o��6[�?�}�'�bG  `�j��Wk�b蝲�1���+�!v  �4����z:V�  �z� �I��m�)%�ߖ��[   pT���ce�c�Qw���:����   ���k�:+���f�r�L�H
��   �j.�(��t��y�  ��a�  &��k�\��ߒ�9v   ��AIK�c7��H�����[�bG  `�5����$�BO�K2��fz��ٱ�   p�I����|+v  �k1p  �N�ҵKM�5IU�[   p�:ݵU��r�R��;;>=;
   ǡmCҒu���l���l��ߑT�� ��2����L!��f�p��LLvӚ4s��Us�2�X�����h_���{����!   ���  L"nMK���I�E��  P�J���i�e�5�m�]����۳�a   ո��$�\Z$�%��+�:v `zI�)I���`JB82NO��8=��瘤p��L��� ��Q{����e����fGF����R�*����Uʲ߼���,S���>0�\Z_S]u�_�q(v  ��p  L��pw����W$�h�   L�~I��|�����oݽ��m��   ����uu9�Γ�%r-6ӻ%͉� (fR.%IP.�W�����z���=��|��NTǨb)S1�T,�)��_�u���X�8-���#+��]�\�;  �{   ���UM��#�ݱ[   0i�ۿ��O%�txd��}��Ծ�Q   SY��>_�U�o�w��wL�H��bw ����M�$�'A��G�|?�>=��f)�I5\L5RL5t�-�w���<W�l����!  `zc�  �jn��mn�?J:3v   &�Nwm5�&m�\��ӱrw�(  �ɨᣫf&#�;��ȃ-�k���$%��  �K0S>��咠|��%ʽ�����z�d��0R�4\,ih$��HI�#%������U�ׯ�Q�  0}q�  DӸ�K�,��dͱ[   0euJ�f��n�J�u�ƕ�%�)Y  0m���g��s_3f?[���4̔��'����dt̞O�sA	�uHr������)ip����"���됙-�w�wb�  ��{)   ��ew~��p����[   Pv�Kz��[�����}R��Y�0  �ո��$�\Zd�.-�� v `�|��o��9q��J��[N[ǉ�2�P������h`�����t��le��+��  ��f  ���s��-��H��n  ��q@����gf��[x�nq��߿}8v  �Q]ޞkij9ӕ�'��]~�d�Kj�� ?fR>�9u��O��/<�t �,s��th�ݻ�    IDAT�������F8���d�W���)v  �^� �	5g��?����!   ����3A��\�P�'T
�wm\�d<=  &�춵'%�s��2;W�Εi��B�6 ��yy�^ȅߌ�_�>�=�0^�ԑf��������R^<��}�{A�J^!  L�e  `�4-]�g&�U�   �M4�i7mw׶ ��I���|�+v  ��?��ZU��/4��k����dͱ�  '�L�%��r��_�z��+w��PQ������{Y�{�g����c�  ����  L �9K���H���%   �[eR�K�M�Un�2���P�g���| v  �d.o�5Ϟs�_��"�-pi���%�n�)(	����_���Q;�Q���������e��w}����텯�8�  �7�  `|�mH���.����)   �8(�􌹞4�Sn�� =9�K�����Ď  �k^���UqV��r�9nv��Βt����} �c�S!��"�(��'A�|2:^��u�-K3׾C���?���R��	��U\���?9�  �/�  `�ܴ.߼����li�   `��|�L�ܵ#ȷ+�m]�u���v^� �)���5������m����Od?KR9 �&���8i�ho��0�ճP��N���i�W������!  �<q  ���n��rp`��]�P�   `��7�)7=e�oϤ����j���g�;�� ��������tN��� ���96��>v ����������|�p�:0�����?���!�Ǯ��ʆ�+TΔɶ&I����Y��	  ��  `̝v�ݕ���L��   �BRI/��K7=�rNY�\�l{Aw-/� `�kې�${Nv�oW��fo���n:Ǥ�%�c' ~[L�|��\�B>yՠ�"�(	L��h�����C�)ĳ��C��\�BU����\.� #w  0ָ�  ��¶�n�n4��n   ʉI}.m�i��vȴ�3�H�<�ױ|�>  &��m
�Y�<%�/�|��K�7�ΑT9 �
I0�s��i�Gy�O��ePֆFRu��ׁ���)x^T64�0#w  0��  ��v    ��$�8r;<�W�]�u����,r"  c���5����[���b��:MR�� �����$(�U�GOa/��s��`�����ۯ�b;�#�//��I���Y��\�,a�  �
w  0&N�rU����>�}0v   �W9$�s2�0��]��.�hn/fI�W�g���  0�4��nI�Nβ0ϔ���N1��=���f�n H�L�\���[N_p<ܥ�}�Գ@�k�j���G��<���T�Kf?��%/}��=q�  @9�$  8a�6z��C҇c�    8nEI�&풴C��L�K��i����w�����2 `L�v�ݕ�[�h������#'�K��N�4#r& @����_q�zE>Q����\��|;@�.���9�}�҈���G�MF�  `�1p  '�u��}�F����   `��K����^���,�Up������������"7 &��n��r�P��,I�Y�S]:�d���3;���\���	 �S!��"��p��z� �'�\/���ރC�S ): /���?GF��g##C���O훸:  Pn�7
  ޺��д}�7LZ;   @tC��Lڕ�:-h��;�՗ۥ�;Cf��f'/���ر ��3��UŬrn�U���[e6�M���>������-��' �4��|N�|�B.(����|d��`
�=0�]{�弶\Ti��or�~R��z����˗�t�쟘:  Pn��
  �"�9K׬�ly�    S�I}.u�� ^��L���;�m��Yg)�}��o플��`��v�ݕ�C�J���y���y�I����Ms�:YR>v/ ��^>����Se>9<fOT�O8�@��,ꅮ�J3&��Ӣ��=���GF��f�?���o�:  P��7  ޒ9K�~N�?��   ����k�I{M��f{\��2��=A�׃�����|޳[-{ձ�M���s��w�	����fg�}�)kp�l�$k��l3�vi��FI3bw �]0Se!���÷ÃvF� �������ܯb��N�v��C�������T���d���Z�  ǋ{�  �5/]�����    �:�IꕴW�=2�k�W���{C�=�|o�'-%�ܭߒ�A^6@l�W��Ns�����>ە5��l�7��`�l�7H6[R�F�<� e�c�ꊜ*�9��憋��۵���K�J��q}���}�L��kÊ��*}  �xp�  �9׮�En�cw    �8��'Ӡ|�}w�Ӡ��̽ϥ>s�I6����՗��\6�˲�R������mK��_ SҼ�/T�WV泴*W��4X}0�gf�&��L�n�7Y��UnV���ToR�KU��5:T���� ���OTS�WMe�1; ����T�u�S����I��%?�?o�U)T�����w�m�  �w� �1kn[s���.)�n   �)����2;$WѤ�L�L�/I&�IRf:`R*�C&q������((�^��,�3�\!;����>��l8ͧCŐ�6`�������3�(Kuׯ���
E��U��,�,�*	�d�,IrY��I3B���U�Y��*�T���j�f&�W�LA���.U�T)W����7  �[!����pd�^��; ��ᒞ۵O�s(���lt��Y�Z�r�L��]n��ǰ  �1�  ���,]��L���
�[     'lĤCG�����[�xwi`��P��U������f�Q��p�Rz�� `
	f��̫�����U��I 0������bg�=�J�������Z�B��tcφ[�f��  @c�  �T�5w.�$<�/�        �De!�����TU��xv ��K{�ջ��^�c�Ӣ��='�}Be�,_U���+��� �2�]h  �������ǒN��       �de&ͨ,pJ; L�,s=�R���i씲5VwI
U�d�ʃ�}=�W<:&�  �%�  �u5|t��\1���w�n       `�yy�^7�Bu��;	 ���ᢞݵO�Kʓg%e�z�軙BU�,W�LJ�{:��Wc� @�a�  ��u�9�Jߕ�wc�        0�̨�k֌JF� 0I���מ��3����%)(�4H!�d������1��  �LpO  ՜��W�       0�"����Fg�ܠ�ϝ�ٵ���`�h��V8�s<ؘ���)�yvN�F�[ض�0�   e ;   L>MK���\��       @LI0��V�~F��+�s  �#�5�U��o vJ��q��\�*�SR�𾞰g����"  `*Kb  �ɥi�>h�/�Wz       LSU9�4�蔦Z��T(��u ��*9�90$�Rn��#����z&OK
��w�X����}�'c  0U��<  ����/-�,�����[        �H�FOko��Tu/� Sѯ{���P쌲���H�����|�B�����������  �)��;  �$�^������5?v        %�j�Y��3���B��l`��g^�;�줇�HYqܾ��)+T4��vݻ�q�  �2B�   0	ܴ.����3n       LU9��T�sN��9���@���+�c5�l|�L����p���CK۪�q�  ���  h���.���       ��V[U�魳t�I�j����k��RWS;��XH����~yVz[j�{uy{n�/  &5�  LsMmko���;        O�U�q�,͟[���|� �8��*�N(?�|���L�@�̳�ϙ��_'��  `�^  &��k�\,��3       �L��T��晚3�Z��@�K��g�`��⩼4<��%�|�{j���Cۿ��	�(  ��x�5  ��9�}�Yi����n       `��V��P��
Nk���/��p1��Q6<-*�3a׳�������{W<1a  ��D�~  �l.o�YZ��q;       ��TW�����4n�v ���
��	e��ľ���ˋC5.���m]݄^  L
�4 �44gN�_����        ��B>QkC��j*b�  "��8�sLY�y6a�̆�+��|����#���]  D7���  D7g随H�ג,v        '*����F�4ժ��3�  �p)�����e�KÒ�|��|�Y�64����'��   *�m  L#M�|�K���jc�        p�f�Th��*pR/ ��֯���(+��yq`�/�T(��O3�z;ny`�  @�� `�8��U��z1n       Lq���No��S�g2n ��$p��X�$��鰲�CI0}���u�q"  �D�>  �����J~A�        ު`����yR�j*#�  �^0�c.��]���FN*�ҿ����  LI�   0���|���Zw�       SҌ����R���
�[ ��R�i����e�,�G$y��{:�P�:cƹ��?��{?�  &'� P��hռ`�1n       LA�L�j����T��7 ��K�8#첗��]�S�����5_���x!  `"0p ��]ޞ��r�H�; ����;��,����;�n��K/3==��R\d-�,QR$[�I۲�CJP,[�DQrl�p;�3�_�9�a�A����ț ��+��Erv���޵޺�9'/zHΐ�TwW���{�h�@�C9Uu�{   �v�tZ��=˱:?�:�1p?Y��6��G��mUU�O��YL 'w c뛛OFď��     �ۑe�Wf�3��p�܏G�{DT�ݨ���Y�[ ��c� cj�3O�����     p;ڭF<tf96�f"�R� PG��0u�X���	QlEV���x��_N� w C����g�����p�    ��X���#g�c��L�@��E��e��ܫ"ʃ툪z�̅gΥ� ���; ���?����Sw     �adYęչ8�����v �N��c�5;�""�D5�.��œO������ ��槟�dVů��     ��h5�x��r�/N�N`���ckT���NT��'7����S�  G�� �ș�>�VE��Sw     �a�N�⑳�1�i�N`L�t���Z�hEd�29+��nE����|���S�  GgT��  ���(���S�;     ��,�OŃ�����kk ���~/u����s�=�A���NUV��/|��: 8� ��X����BD���;     ���Z��s��e�K '�A��Aꌱ�5Gh�U7�r��+ٕ��� 8 �X��ԩ<˞�"�S�     ��ɳ,�m����h� ������3�_UF�{9u��e�ḫ˼������}� ��� c ��)�v     FY#��Ӌ�� ������A�ɐ��vꊷ��({;ͼ��i��3��9 ��1p��[��ӟ�,~!u     ��V#�N/�씽 �����eꌉ�5G�k�`?�����7ʿ�� �;Y�  �Ν�s_\���Dd��[     ���[�x��btZ��) �������z=ʪJ�29�"��+�+�Wֈ��Z/����x�sϥ� �� Pc�v���    U�V#:�d����������7"��߫*���vʬ�'�䓶q PS��@M�?񥟍*~%u     ��v��^�Vӯ�8>�vb{��:c"�ͩ�	���EU~d����L� ܙ,u  p��>�{��T�?FĹ�-     �ݾ5no�p���a<���(J�ۓ��(v�D���?kDcvm���_�7^I� �O ����ޓa�    �j5�x�Ԣq; �jX��ҥm����<��N]�Ϊ"����0+�a� ��y�  5���ӏG9u     |�f#�O/E��H��+�*^���A�:e�孩�	���GU��槟�d� ���@�TYT�#���     �*ϲ��Ԃq; Ǫ,�x��V�R�Y�Y�wQEy�Ud_����?�� 8<w ���O��_�"~<u     �U�Eܷ�3�Y 8>ߺܾ�5nY���}D����se�o�N oT?> |�{.���~��jD��n    ��:�6kө3 c�a/^ڊno�:��R{Qvo��xy4�V��<����[�� x.�@M�����     �����v ��~o_�q��ʚ����:�=�Q춋*�݈�AX ��Q�� x��_�������<�f�G#Ͼ�����Y    �6sӭ�w}!2O�8&W������(J�'iUQ�SW��rY�u���������?H� �7� `�=�d���ƿ��L�^�e1�n�T��V#��<��F��y�y���h7�h6�h�ydYD����������UTQEQT�����3��c0,�7(bX�'��   �I�j�����h6�8��7��ͫ;��?£i��,�ػ�����ḫ\��G�����v� ��5S  �m�+��Yd��0�ڭF�M�b�ӌ���?S�fLw��i�˒n��h��_bn���������� �{����c�7���A���   �ۗgY��\4n�X\�9����𩓼��D��%�F��n6���""�v� �ݹ� #l��SsY��QD�I����g1;Պ��v�O�cn����h5��˻��b�`7w{��ߋ�=�w    ��=��:?�:�1�����vc�`�:�;P���L��>�ḫ���co���|)u ��\p��g�ߪ���DeY��T+g;�<73혝z���u�ȳX�i��L;"�#�ֵ���^�����^/���QVU�P    F��lǸ�#��q��^\�9H��]Ț���Q�S�Ceow*��^D<�� xg.���ڼ���s�p�y�3�X����ܭQ�8\f?JeY�ͽ^\�����.�   L�V#�G�Y�f�34 �^Xƕ����}��Θ({�Q�wSg��|f5����+_���� �^� 0�6>����/��q4�i���L�/N��\'�̷ŷ��ƕ�ݸ��7w{8   L�N/��t;u 5w�/���~��=�f3U��y+3����� �|�L� ��% ���O?��DT�&|��#�l䱺0��ӱ�8�V#u��e\���_��   `̭-N��չ� ��N�W�����O��1*�7���x_��bDk�׮|�7�i� ��� `�T�槟�wU��S�@��[��\����X��J�3z�".^ߋ7���N׃i   �q�n5�ѳˑ�~����˸�s�w�?(R�p�������/ˣ1�~1������7�R�  ��L  ��槿��*2�v��fK3qjy6V��OZ�Ո�q~s!�q��^�vm��j   �1p�ڜq; �V�Ul�����A�v�s8aY���"��k_�Q�wO7��߉��6u ��@ �(��gZ7��"��)P��wF�F����tc?^��7�z�s    �K���os!u #nX���ߏ�^�t�QU��H�t�<�J�qY4fWw���Х���S�  ��� #d�F����a,̴㞵�8�2��FV�eqje6N����~?^��o\ߋ��T   ��,�ӫs�3 AU��c�ۏ�� v�����5�ۉ���)��7�M-�͈���5 �-�@ 0"�/<5�e��#�T�U�F�W�➵���j�����E�vu7^���A�:   ��pfu.��Sg 0"z�"v��ߏ�n�A�S�ۍ���:�P���~#ڏ]���!u ��; ��,��zDe��`i�������Ld��h�]�و�O-�}��՝x�Ҷ�;   �j���`�0����no��A����0�A1�׸%yk:��^D��!��^��i���R�  .��H8��gֆE�|D,�n�Q�ek�q���X����UU�_ۋ�/ތ��;   ��8���s��L������3f���q���b�ݭ������O���h}�ʳ����n�I�; ������̸"��gqje6��X�٩V�N@�eqvm.ά��   ���vӸ`UUDoP��`�~�a�E��E���_�<7�    IDAT٦~��lm�eo'oή���S� ��s� [��?:����#b*u��n5⾍��gm>��<u	�e/_ގ�؊��0    ��O-��L;u w`X���1������c0,S�1����E?uơ�SK�Ο���o���[ `��� ��U�o�q;������b�[��<��K"�<��O-ƙչx���x��n8   prf�Z�� #�,��U��m�6f�����۳Qv�1p/{;�hN������[ `�Y@B+�y��f�}="�畉�j�qn}!��\��a;�ag�_������K�   08���� ǡ,�(�*��֟���(�w��o�{�)uV�]�(�3%�Z��L�ؕ���� &�� �P���V�3aZ�<��\�s����L;��#���{��nDoP�N   [S�q;0V�5/�����[���u@^|���|�q�w�΋��*�����?��n��:��$��3Ql��8������߉��I� �ʢ 9s�sì�Z�3!y�6���B4y�j�(���k7�WvR�    ��{��ce~*u�����uɼ��E��ͫ�e��ۮ����[����ؽQ�㐑+� ��� ��0���̸����8�޻�m�~rwy�ݻ��g�W���A=^e	   P�F�s������9N��7�g�a�a���X�-��=U�G�n]q����ө[ `�� 	�y����=�����v<z�J,��,G�,�x���x��׺   ��+���4�:3U���������[#v�xaBT�+�Q�.9���ў��+_���� &�� ��0/�����_�f�Z�s�Scy���g����\|�嫱��O�   P[y��ʼ������h�[�ް������ ""�<��tT���%�R���њ���n�I�; ���O�md��z;c(�"�m,ă�����V��SUU|�������)    ��4ۉ�6Rg #lX���o���"E�C؁ë�(v�DD=�Ƒw"k�����~�ߦn�I�; ��FV�NDf��ؙ�n��[������eY��]��������FP�N   ��e�ہ�����������K���%v�dyd�����%�R���ў���[ `�8�	 'h񗾴���1���J�eq��Ÿ��Bd�o/I�?,�?�t-�m���(   @j�F��[��`rTխg��A�a������'�*�Q�]M�qh��b��;z�_��WR� ��p� NPg��vDe���X���έ��T+u
|[�و�=��\މ��v�/c    ���\Ǹ��;���8���dy3�щ(z�S���f���_����� &�� pB�|��t�RD��n���l�����gm.u
������/^�ޠH�   0��g9��n�A��2�Et��[\dFXU��ܿ�:���A�9������+�[ `xJ 'd0S�ZV�S���x��Z�t|+��[���}����^�[{��   p�ڭ�q;��`X~{ľ������C@�d�vD�Q�S�J��k[�5"�Z� �.��I�ē͍���G���)p��,⾍�x��r��mUU�s�\�ׯ�N   )k��qv՛aTUU��"{�7���0Jgف1P���L�qh���~kj����߸�� Ɲ���	����L�ScS�f|��Z,�uR��ɲ,>x�j�O��k�]�J^   �7-�x����"z�"�{��ڍفq�5�"�fD9L�r(�`ofؚ����oR� ��s� N�慧�]�e?������L|��j4y�8W���/^�aQ�N   H��g����"�[c8qUq0�5`�w��`ՠ��V�C˧W�v�o>�׺�[ `��� ���g��DYV���N#���V���l�8Rk�񃏞���rt{��   p����pB���W��{��;DQ�d����NDU��D�`m�X������- 0�����e�WR7��j7�#���L;u
�٩V�ࣧ���r�t��s    ����GUEt���;�Θ}0��p��e��f���9�jxU9�;�?��|R	 �����1:���ϗe���h�n��Z[���_�f#O��nX����_�����)    '���]�N��k�[�a{o������2y8���b�jD���@Yk&�ş���o��[ `\�� Ǩ(����S#�7��˩3��4y��Û�^��o��   81�Fn�w�7(b���A{o�a�$�z���ZSQ��jЍ�3�W#�� ��� pL�>�{��T�ՈXL�������Vc}i&u
$��+�⵫�x�%   ��Z����ͅ�0�*���y�}����0P+e��Ո��+0��|��Ǯ>��?J� ��w 8&��ޯU�q;�o�ӌ�>��S��)��έF���˗�S�    ;�᝕e��a��c�;�noeU��%@��ȚSQ��K���g����#⯤n�q�; �'��7���ZD<�:���l'>��z��^E���oƋol��    8V�]����;|�B�n�֠}�``��HU�ܿ�:�����as����_,�s� ���n�\�q;#mci&>t~-��g�:�a�   ��,��n�3��*b�wk�n�0Z�F+�ю(��S���ϵ�S��0u �w 8eY�Ff3�;���޳�:F�Cg����x��v�   �#�n6�3l&IoP��� v�����GQ����=e��(Q��ET_��|q�#� ���<uo��^��F��nY��=+q��|�����z=^���:   �H-�v���B�86â�݃A�9h��I ܆b�jD9L�q(Ys*bj�W������ Ɖ� p�e��a��ʳ,>|�Z�/ͤN����{W""��  ���iy��x�����A�toڻ�z�"xgyk&�^=޲[{�W��"�� ��� p�>�dscc��8�:ު�g���cma:u
��W^��_�M�   p$�]������pW�E���o_i/�*u G���ػQ����~3���ҿ��˩S `\�� Gh}}�φq;#��g�7��
���[�aQ����S    ��T�w��_��~/����w0H��qɲ�Z3Q�kr|��m�ss1"�^� y�  'Y�K� o�j���7���|��Z,�vRg    ܵN�4�,����ūWv⹗��}�z\��g�0��LDd�3�*"��'����#�* ��'�y0��'Sw���y|���X4ȅ#���6�٩V�   �;�gY4�ŘHEY�ͽ^�re'���x��v\�9�AQ�N�$eyd����7����� 0.|4 �JU|.j�r�]�Ոxx��X���Gڈ��ވ��H�   pۚM7�=â���~l��b�ۏ�J]�(��3Q��3�D���G���� Ɓ �O<����x5"N�N�V#��?��3��)0�v����R]�   jf�ӊ��.�΀˸�׋��^�R� 0���ke=�Nd�a֞��ʳ��F� �;��#����sa��h6���q;���v<~~-2   j��;	e�w��7��_��_�5n�=���	�V��,�_J� ��� 8U1u4�,>��z,�ÉX_��O�v   �K��WĜ�������+Wv⹗�ūWvb{�U���:�ZSYM���(��_K� ���A �Kg��W�����*&�<���\�����)0q��ū�ƍ��    �rjy66��s	������v7��zQ��� ܹ��U���ɚSSK?p����?�[ �Κ� ����W�2n'�,����k����[��� ����S    �W����񩪈��^\�>����e ��5EM�հ�j�"�� �BM�� ����WS70�>x�Zl,����y~`=ZM?^   �/�o��eW���\��/m�p��ƭ��PE9�}����B'u	 ԙ ܅�'�������L�O/����0�������1   0�2�/8BeY����^�ׯ�Ơ(S'0��V}�f]{�[�O�� �:3p��Ш�_M���:�:�^L��ii��YJ�   �|@��rs�_����x}/��� ��َ��3�D�)u ԙ�; ܩ_�UE|6u�ii�8��:�.�7b}�>D   ��c������k�݈�/m�`h��I��v����/<u*u ԕ�; ܡ���D�Z�&��T+>���W	È��}k�i��   0q\p�Ne�^ى�/ތno�:�	��j��mD��; �����Y�z;'����#nD���8U�f��54    �ƍ�^|���q}� u
 �,oD4ک+�*�v9u ԕe ܁��Ϧ"�O��`��Y}p#f:��)��X���N-��    �eU�N�F�E/]ڎW.oǰ(S� @���ǰ���/<�P� �#w �{������L�G�Y���N���8�+�S�3    ަ,�9��n?������K� ߖ��"�zLުa/�j��� p��� FL�B9QgV�������mz��Z�~�   F����x}/^��W�9Ydͺ��~9u ԑ� ܦ�_��BD���L���v<v�J��tZ�x�  ��;�?,��ߌ�7�S� ���Zө�����>�� ��� nSc��ň��G©�V#��p=�<K�ܡ�+���4�:    "\p���t��o^��� u
 ���ъț�3��E\q��e� �)�곩�Y���k1ݮ���]=vn%Z?~   �.���lu��7�����Ț��IW{�Q�h ��� né_X��O��`2�j1���z=�ݵ����{WRg    DP�N`�TU�k�v��k��? u���3p���{6�x��Rw @���m��柉�9v3�x��R���Z������   ����󦢬�K[qu��: n[�7#�V��)�Q>u ԉ�; ܆�
?tr�y�=up>pn5ZM?�   ��e�F@oP��_�����) pǲf'u¡�E�B� ��
 8���,F�O��`�}߽+1�� G�f��]N�   L�����'�~o�x��k� �^֚J�ph��ྍ'~��Sw @]��!����N��x�X��3�s�3�ctfu.�����   ?��a���⅋[1,|�����fD�J�q8� �����3 �.����|� �[�Ո�[M�����]�,K]   L���'��^/^x�fe�: �Lͮ�� �!��!���33�3�;o��_�Vӷg0	f�Zq��B�   `B�R'p�n������Qٶ0f�f��E���_z4u ԁ �`�����I���:�6+��y�ܽ��,E��H�   L ��ru���0��FD�L]q8E?�j�; ��; F��:���n5⑳˩3���3��   ���e�N�������� p��f'u¡UÞ�; ��; ��^�r;��������]�f÷e0�N��z{   ��+���ҍ�x��^� 8vY�>�(]��/ܓ: F�% ���������������X�I�$��=+�e�+   �Ic�>ޮlu���Y�u��U�^�l6�t� u��� 	�?�����l��ع��@bsӭ8�2�:   �0;]�que��_�M� '(���NqHU���O�� �Qg� �#��9�]�N��:�Y�F�;   pr��8��38b�� L���I�px��'�|�����`� �a��*N���Y���=k.6�tZ�8���:   �0[{��	!�v &Y֨���j؟�w?�� F��; ��<��t��ӣ���N F�����   �	�i�>6���xy#"o��8�2��}*u �2w xUT?����sfu.f�sA 8�<��7Sg    �?��~�:��t}��� ""k��w��p��U�� F��; ���_��B�;/�<���,�� FԽ�s1ө�u   `l��^k7v{�ͫ;�3 `$d��ܣ�����J� ��� �Ec��Saeȑ���btZ����ʲ,8�;   pr�mw��RWp'��z��m� �MY�F��/���I� ��� �E�ϥn`�L��q��B�`ĝ^�u�   81��������nw�\�1n����>�c)��ϧn �Qe� �*�����G�.G�g�3�����    '���~�n�~o/���u; |�z]q/?�|����w`� �`����I���X�����L��&ά��t��:   ���0��38���0^�h� �&k�S'Z5�7[1��� 0����T�O�N`�<xz)uP3�o:�   ��+[��	��n/��Ei� �Q�Be���Ϧ� �Qd� 2w���l'V�Rg 5sv�w   ��l��\qa�A/^܊aQ�N����͈�F��r�S� `��9 ��^�r;�������κ�ܙ�   '��k{�x�a�_��v 8�����Ъr���t� 5� �]�Ƶ���������X�s��3gWg��j��    &�~o7v{�3x�aQ�o�`h� ��5�3p�r�p�'Sg ��1p�?�:����i�ہ;�eYܻ>�:   � ��FYV�3�[���/nEoP�N�Z���	��,����w�2w����t,�uRg 5w��|4�,u   0!�2�luSgL�aQ�ol�A�: �'���=��'��� ��� �����j�����N-�N �@����չ�   ��ts/����e/��ݞ� p'���9T��S����� �Qb� o�of?�>rg;��G澍����   ����x��v�e�:e�e/\܊�� u
 �XV�+�UE��gRg �(1�������������12�i���t�   `��E\���:c��e/�a� G!���="�b��� 0J��-�*7p�Mw���4�:3�6|p   8YW�����ΘEY�ol�ށq; �F��Q?�x�f� p|��M�\�'+�SwP�֍P���2?����   ��y��N�eꌱV�U�pѸ �R�5R'ܖ�̞Z_�X� � �~���𵑻�j�qvm.u0���   8i���.ތ��R���aQ��o�~ϸ �T^��{DŠ�S�+ `T�����O�@��]��F��� �ԙU�   N^oP�K����q?R�a�_܊no�: �NV��{DY>�� F��; �)�ܹ;Yqnc!u0�y�˳�3   �	��īWwRg��ޠ�o\�}�v 8Yu��eU�#q���[��1��Wq 8&��Y�,>���z[[��N���x�]�K�    L�;�ƍ��������oFP�N��V�+�U1�_o\�[ �0p���h�埈�z�t��9�6�:� Ks���n��    &ԥ��ڵ����w0�.nŠ(S� ���j6p�(#���T�
 � UT?���zk���8�:�g\q   ��ՍW��DU�.��k;��ś14n����oW�?�� FA����q��M�@�ݳfl
��3+s�gY�   `���9��/o�BUE\�����  8Y5�W���#*�`���8 ��~���죩;��,sM8Y�fK3�3   �	��׋��r��=e/]ڊ�7�S� ���j8p�r����?~ u �Vï� p�v���������tL���3�	sj��   Ho�ۏ��v#�{��)#�7(��ߌ��~� �Ly�qUU���x5�* G�*㏧n��κ�$��8���   ���2���MW��bk��x�f�S `r��{DTÁ�; ��_��(eُ�N����<��Sg (˲X_r�   Uq��^�ti;��J��LUE�vm7^��âL� ����j�é  �z~���C����t�y�:�P�WfS'    ���^/����q}� uʉ������o�խn�  "��ܣ*[��׈0�j�U �ƙφ��}    IDAT����I�A}m��$�2?�V#u   ���2^��/���A�:��UUĥ����nD�7L� |[M���F��� ����hE$u��l䱶8�:�p�ˮ�   �i{��������(�*uα���k�݈7n�E5�������#������ �R3u  �T���d�8s���#��C`<�^��W.o��    xGUqe��wbmq:�g�����jX���qs��: xOyD��#n[�c} L4w &ZVV?\׷������(X�i�T�}��   FWQVq��~\�����T�-�D�Y���2.�܏k�]���,��_���R' @J�{b  G�ןiEߟ:�zj5�X[�J���(   PEYŕ�n|��k�ҥ�����b(��ڵ���W���-�v �����r�z�3O�O� �����Z�.�e����td����hX_��W���    8��������^/Z�<��:�8ۉ٩V괷������Al������SQt0"^J� )�0����g�ܩ�ג�ѱ2߉f#�aQ�N   �m���+[ݸ�ՍV#���v�ϴcn����_]��ck�7vb0�� H�*?_N� )�0��*>���zʲ�����ёeY�.Lť��S    �ʠ(���A\�9����v3f:͘�j�t�S�F��Ѿ]�7(b�7��n?v��1pD  �G���]6 L,w &V���(KB3�h7�3 �f}q��   ;�a���GD��yL���j��n6��̣�g�l��Y�o��,�*"�����"�����������^��n�x �H���G"�,"�rz &��; ��ןie7��Π���S' |����Ȳ��#N   `��e��� @-���]Y,m^���K�Ƌ�S ��  �����J�A=�.��0z��<g;�3      8U��J] )�0���x��e@
�0o�      ��,�����(�X� H����TUa��Y[4F�ʼ7L      |KUU��NU�6 0���TK@=-���kq����      �AUUN�  )X> 0y.|���Π���:� ޓ�O     ��r����M� '�����W�����O����T+u�{Z��N�      0"��w�*#�|4u �4w &N��WxqG\E�`ua*u      G�����8� L���>���z2p�`v��V#u      G �
 &��; ���]p�,����:�;     @TUꂻW���N ��f����]p��eY�⌁;PKs�      c0p�x衟��_V0Q��(k�����������L'�<K�p(K�8     0ܫack&>�: N��; %��+en��L;u���M�����     0��`�1��h� 8I L���p��i~����     &�8\p���[ &��; ���>�:�z��j�N �-K���	      ����=�����b��D���`��in����E�    �I6&��#"���R' �I2p`�dY|_��g�ӌf÷M@�,ι�     L���WUqj�S�7�� N�� c������8������r���v�ӝf�     �$���dI�����{j�@��,���n��
_Co}����+_����޵7��>��Z�@�#Hb P�5�|��>/(ɢMR@!3��/�'��!��"DdU�?ߓs*�0?�o�+� lw 6Ƶk�\o�J���W:�J^��     ��j�G��t��� �,� l����;Wr뺁(������/     `C�\�`���w���a����ڊ��n`=ݼ�S:�Jn]�-�      PFm�G� �� l����q%7܁5u��     �fʕ�sJ[� �������63W���;�~d�Ӎ��     �)��s�s�Q��/\g`#X: ��ۿ�����t��ƞ���v��n�     ���{i��^�{ `#��^9��D��O���v��gr��^�     ��l����?/�  �`��F��iV���t��E ��yw     `�
�]��c� Xw 6B��ߔn`=����[�}Q     �@�/]0wMJ?-�  �`���h~R���tso�t�3�q͟c     ����{���� �� l�l�Ε\3p�ܵ����jJg      ,ON�KW�]��K7 �2��ܹ��?.��w     `��
���ѷ����^� X4�- ���؉�+��z������n^�-�      �<�ҁ{�M���t ,�� �{����ADX��Ԛ&b����M�    �M������oJ7 ��Yl����.`=��l�N ��.�     $�z�� ������-w�doǏJ@\p     6J��s�Z� �j��5���+����P��     ��)�NX�&7?*�  �f��hܹ�����	 sq}ןg     ����{?,�  �f�@�r��t��w�M�Į?�     �M���G��N �E�p �~M��t�iJ �ϵ=W�    ��SD������o�ӿ�Z: ������_�����F��Ӗ�;P�k�;�      .�|�=""rL��?*] �d�@�vg���\�֖�;P�k�.�      u�n���P5w �����n`}�����     ��_p�H9��t ,��; Uk"}�t�����ގ�;     �6`�)�B P5w ��#\p�ʶ��T����;     P����	�4����mP�&·�y.������     �r��s��-�  �d� @�w�l�1p�k�     �.����]�)�  �d� @岁;W�#�N ��mw     �r9��=""r~������ �E�p �^���VD�Q:����ہ���     T/u��$mN?v��jY8 P�W��oF�o,se�����_�     ����G��~P� ���z���N`�ٷ���jJ'      ,L�7gྵ�|�t ,��; ��N��K7��rX�u���+      P����޿Q� ź�z����g���;P�]w     �V9G�t��䰉 �Z� T+G|�t�ͼ���VS:     `!�]o��h"�D P-w ����2��w�6[��;     P����� �2p�^�1p癤l�Tƾ     ���]p���� �(� ԫ��<��7p��;     P��o��=7��� �(� T+G��L�>�N ����     �UjK,U��7~�_���� �� T*7MxϦ7p*�e�     �(����,��� �E0p�Jo���x%"�Jw�޺�qo� �۲p     *���tByk��� �� T�O�[�X]�K' �U�     @}rjK'��$w �d�@�R�^:����.�ui��    �m��H���	 �� T)5�j��_�܁�d�      *���S��J7 �"�P��I�<��#�d
�#Y�     ��9"m��&�R: ���:�������}���1p     j����?�]p�J� T��-e�df�T$y*     P��o��=7� T���*��w�c�����T:     `���tA19��� �� �)��;s1u��Hk�     T&���	�dw �d�@�\pgN\pj�u�     @Er�ț��n��; U2p�NM~�tup��E�9�d�     �#�]�Ҟ��?���# `���Sܙ���;P�I�GΥ+      �'��tBq����� 0o� T��N~�tu�u�u��|a     �K�f���ى�J7 ���P�q�x�t��6��v@%��H     ���h������P��ԿX��z��>Rʥ3 ��x�^     �9u��s�m$ ���; �I��~yc�\qj0���     �H�ODDΎ Pw ����F��b��`4�&/     P���J'���F���P������\�����N�    �z����s�� 0o� T'�-��b�&.�kn2��R�     ���)"��+V��� `���N�p����k�b4-�      07�s��O�H6 T����lm���O܁�v>4p     �{�?I9�H Pw ��s�b��b�����7y    �z�-��J^(  �f�@��Nf��>Ŵ�Kg \��;     P��#����4.�P!w ꓳ���p�`='mt}*�     0��Qn��K7 ���P��㷘��؛$�z:NK'      �M�=�������; ���7�n85p���ț�     @=ܿ�i�f� �7w ���s���`�M`=�\�K'      �I����%���_�P/l �����N\p��p��x�M^     ���""��X5�kp����P#w��R̺�t�S9v�     �H�=y�����K7 �<�P#�Lf!cW܁�r|n�     �#w��	+��M�J7 �<�P�����ۥ;����5 `}���l�M^     �9G�}���.�Pw �2�u������X#'�H9��      ����"�g_�I[� T�������~ica�G.!���b\:     `nr��گ���	 0O� T�iw�Y�񴋮O�3 ��ѹ�;     P�ܷ�V�V�Pw ���7K7P���t�_ur1�Yۗ�      ���"���W�� �����4͖�,���c�շ:(�      07��9��I�7p�*� T�I��,���w`�����|\:     `nr�sگ��� ���; ��7JP��7N��vp6��O�3      �&�>��:M�� `���J�f�tu�̺���� _��ɠt     ����Ed��~��V���P�&ǵ���l0)� �m��     T$w��	+/7�����P�&�_�X��Co� �i�t9��      ����J'��&�� U1p�*9����¹���ώ/K'      �Q����+/���Pw ��le���p�qm�Jg |���(�Ӯt     ��䮍���5Mv����P���_�X
W܁Us���v     �.���NXM�N �y2p�*M4�,���t��'m<���     �.�����
O��*� T%��,�!)�J�\�N      ���G��t�zHa+@U����,��x]�Jg Dۥxt:,�     0W���'�� ���; UI�[,G�'�P����2RΥ3      �*w��	k��.�Pw ��;�t|1.� l��r�;�,�     0_9E�m銵��q���P�&�N`s��}v<�Yۗ�      ��ϯ�{���y�t ̓�; U��k�3k��] ��9ǝ���      s����'�4[M� �'#@ ���kK�;Pʽ�˘��     T'G�f�#֌� u��@Ur�嵍�2pJH)ǝ���      s��6"R�uc+@U��P��[�,��`}ʥ3�s��2f��     �ݤt���ۥ `�� ���6�*�W܁%J)��C��    �:�nZ:a�8@e��P��k�wx6*� l��    �Z徍�>yZM�4� `�� �J�^�X���q�Kg ��R�yt^:     `!\o�"[	 *���l��n�|]���rR:� ��Ϣ�S�     ��0p��&�J P/l T%ǖ�6�8x<*� Tn8i���e�     ���)"��+�T�]�  ����d�)����X�>{9��      X�۟A�4� `�� �K㵍2�.���tP���Q�\�Kg      ,Lj}�ze9�J P/l �%�V2�����_�9>|pV:     `qr��g�+�V�[v� T� ���p��2FӶt     ���n�t �"� �d��q|1.�Td������      �Z�� ���; ��K' y��it}*�     �89E��� �
1p ��óQ�ɣ�gwx6�óQ�     ����t �b� �(��]q�M�r���t     �¥�� �"w �9{xj�<�>;�iۗ�      X��"�Y�
 `�� ����I�g]�`M=L���t     �¥v\: XA�  p��w�饔�ݻ��3      �"w��	 �
2p X��\_�����M��      ����~V� XA�  0�vq|�qz��;L���E�     ��Hݤt ��� 䳣��	���S���GΥK      �#�� ��3p X��qLf}�`�w�$&��t     �r�>"��+ �e� � 9G<8q��z�N��:,�     �4�s� �j�  ���t�¦m��?-�     �T�5p ���; ���>�F�3�����h�T:     `ir�"R[: Xa�  v��t������K�I     ���z; ��� ,��`��i�`�<L��ó�      K��q� `�� ,�+���̺>~��q�\�     `�r7��}� `�� ,���(FӮt�~��Q�Zo�     ���v �I� ,A��\q�����q6���      X��#w>' �:w �%yx2��K�3�B���q��]     �͔�ID�� ��� ��O9�]�� 
M�x��q�     �bR;.�  �	w �%�wt)����)��?9��w�     �P���g�+ �5a� �Dm��+�Q޽{�co�     ���v �i� ,ٝ���]q��p��Y<z<,�     PT6p ���; ���]��G�3�;<ŧ��Kg      ��YD�Kg  k�� ��;��C�.G�x��q�     ��r;)�  �w ��.ŽCWܡFӶ��||�K,      �#w� ��1p (���Et}*��QJ9~��QL[��     ��4"�L x:�  ��}�{���3�9z��q���3      VBjǥ �5d� P��Ë�u.=C޿�g��      �!���a  ��� ��)n?<+�<�O�����'2      ���� �U� ��d�I[:��ǃ�x�U      �R�y�- p5�  ������������'�3      VJ��/� �)w �pz9����ur1��۟EΥK      VKn}�	 \��; �������	�N�x��A�ɺ     �r��MJW  k�� `E�m�?�,���Yo�>��K�S      VN��J'  k�� `�|��,f]_:�
Ӷ���QLf]�     ��#��� ��3p X!m��g�3�/1����G1��     |��M#��^ ��1p X1Oqz9)����K��b8iK�      ��4s� xv�  +�{��s.�DD�r�u� c�v     �����~Z� ���; �
M۸spQ:6^���b4+�     ��R�z; 0�  +���M�������׷�l��     ��ˑ�Q� ��  +*���;)��O9��ȸ     �I�v�S� ��  +��r�Jg�F����� Ά��      O"�� ̑�; �����M����>�[��ܸ     ����E��� @E� V\�r���q��ެ���?<0n     x
y�z; 0_�  k�l8�;�3�Z���_t�c�E      �XΑ�I�
 �2�  k��g1���3�:�Y��� c     <��M"r*� T�� `M����O�#�\:�1����hj�     ��lX: ���; �����ó�P���4~����̺�)      k'w���s `�� �̝��8:�΀�vz9��nF�{d&     �U�� ,��; ���ݓ�:W��to�>�θ     �Jr�"�i(oZ{    IDAT� �R�  k��S���q�K��Z�t��=�      \]�y�4 �8�  k�|8���΀�q��Y��Ը     �Y�����  *f� ���^����ur��Ν����y�     ����qD�� @�vJ  �l�p�$n�؋���h���K�ۏ�l8-�     P�y�  �X.� ����|����$�_M�x�G��      s��iD�Kg  �3p ��p���?=.�+��ro���i[:     �i6,�  l w �J�\������3���'�����h=�      `nr�F$ǅ ���)  ���?��[7�⻯�*�E|��q�9�(�     P��z; �$�  �y��Iܼ�/?�t
,M�r���Q��K�      �'���i�
 `Cl�  `�r���'G1�x< �a8i����     ,HjG�Kg  �� �Bm����d֗N��:�Ǜ<���:      "�ȭCC ��� Tj����b��S�;�ۏ��S�     �j�v�} ,��; @�F�6~s�0��q�ԣO9~��Q|��qd��     X�i6, lw ��]�f�#[S�ᤍ7?؏óQ�     ���v�=1 X.w ���r���t<���a����1��S      6B�9: ,��; ��8:�;w�Kg�SK)���;w��O�D      ���D$�� ���)  ���#���G��N�'2����O�\m     X�4�N  6��  ���(~��a��6����0����q;     ���n�z; P��; �::��>92rg%�)����w���S�     ���f��	 �3p �PG�����G���;��b4�_��O�i
     PB�ۈ~V: �`�  ��b���0z#wV�������c4��K     �R�lX: �p�  ��ro~��Y_:�5�����g�}�     �����ݤt ��� ����7?؏���l���l�|�a���S      6^��� �g� @DDL�>���Gqz�"��v)޹s���(�>��      ��� +�� �?k�o�>�ǃ�)T��b�����?u     `U��0"r� ��)  �j�9��{'1m���Q:���]�>;5l     X59Enǥ+  "�� �����Y\�����;��ó9�ǻw?��      ���v `�X* ����o�?��-�j���9���>4n     XE9E��� �w  ��h��/�ۏ�'��)����a��w���t
      _!�F�Jg  ��N�   V_�9�p�$Ά����MӔNb���]�w�$N/'�S      �:9E��JW  |��;  O��� ��6~��W�ƞ%���s|��">}t)��9      �i6���Uc� �S9N�_�}?}����ϗ�aE���N��)      <��"�ƥ+  �?�  <�>����8���������]:�B�m���ÓA�      ���� ��2p ��N.���>����[/?W:�%J)ǽ�����yt�7>     �JN�g��  _�� �g��)޾s����w_�ݝ��I,���Q|��qLf]�      � M�Kg  |)w  �b�t�����_���|�`0n��'q6��N     �R���  �J�  �Mۧ����?��}��x��^�$�`�����Y<<Dv�     `���0\o V��;  sw1�ś���܊�}����jJ'q]���G�q��2��MN     ���z; �� X��#��|�����/?W:�'�R�{Gq��E�}*�     ���� \o V��;  5k�x��q�98��~��x�ś�������YL۾t
      s�S����  ��� X�����~r�x�Z����篗N�r����(>�?�Ѵ-�     ���0\o ց�;  Ku>�Ư?:�o]��y�x�ֵ�I+�O�.�     T.�.r�z; �� (�l0�_}�(^y�F��/��D)�|w.bf�     P=���ub� @Q'�8���7��{�=o��\4MS:�J���ώq��"�.��     `	>��>.� ��� X	��Y�{�$n���^}>���󱻳U:�
�q��.b�d)��     �I�tP: �� �Rfm�ŝ����K��w^�/޺V:k-�����E�^NJ�      P@�g�;� ��� ��ԧO��d��v�[/݌��|���#�יu}<<�gǗ1�v�s      ((�� �!�   V�d�ŝ���{x/޺�y�V������jJ�����q<8���q�\�     ��r7��g�3  ���;  k#�Ǘ�x|9���������x3^}�F\��.��t��Y<z<���aL۾t      +#�� �-w  �R�9N.�qr1���[7v��n�k߸/޺V�nq��6����a'm�      VP��#RW: �J� ��`��`�Ɲ����ݎ�n]���/ݺ���+��L·�8�����0c�v      �FΑf��  Wf� @ufm�Gq�x�[M��ܵ?�޿��^�lo��j�����q�\L��rm�J'     �&�l���  Wf� @������$_N"�<""�v�����x��nܺ��]߉[��bwg��������4����p�J;      W�S�٨t �31p `#��>N�>N/'_��ww��k����{��qmg;���_��?��lE�4O��ק�I�i�Y�I�i��Y�)��      *M��� �z3p ���v)κ��g��&���h�>��?�눈�s�)Gץ�R�l�     �"�>r;.] ��� ��RΑ�ї.     `ӥ�eD�� ����         \]���ݤt �\�        ��ϯ� ���        `M�n��Jg  ̍�;        ��J�A� ��2p        XC�G��t �\�        ���z; P%w        �5��Èܗ�  �;w        �u�S�٨t �B�        ��4DD*� ��         k"�.r;.� �0�         k"O�Kg  ,��;        ���,r7)� �P�         k M.K'  ,��;        ����8"��3  ��        `��H�A� ��0p        Xai6��}� ��0p        XU9E�KW  ,��;        ��J�AD��  Kc�        ��r�"���  Ke�        ���t�t �R�        ����"w��  Kg�        �b��t @�         +$���Ԗ�  (��        `e�HS����e�        �"�l���  ��        ���"O��+  �2p        Xi:��T: �(w        ��r�"���  ��        ����ȥ3  �3p        ((���ݤt �J0p        ((M.K'  �w        �Br;�Hm� ��a� ��a�β9� 
����$�2�}POR�' �*�l��{      (�ї��  �"p        (��KD��  �"p        x���k�
 ���        <Y_^"�W�  8�;        �e�#�k� �C�        <Q�}���� pHw        �'ɶF��z �a	�        ��� �_�        <An׈�U�  84�;        ��e��z ��	�        �/�٪g  ��        ���G���  � p        x���DD�� p
w        �ɾGn��  �!p        x�~�Y= �4�         �m�hK� �S�        <��{;  !p        ��ܮ}�� p:w        �����K� �S�        �Q_/٪g  ���        �^�G.��+  NK�        p'}y��^= ��         ��[�v�^ pjw        �;�˷���  �&p        ��l[�~�� pzw        �/z{o ��         _��-���3  � p        �����T�  ��        ��r�F��z �0�         ��}�� pOw        �O��kD��  C�        |T���R� `8w        ��˷��� pow        �ȾGn��  C�        |@�}��  0,�;        �;�F��z ���         ����  �$p        x��n}�� 04�;        ���v �'�        �A_/٪g  O�        �;���k�
 �)�        ~���٫g  LA�        �+�#�K�
 �i�        ~�//� �Y�         ?�}�ܮ�3  �"p        ��\^""�g  LE�        �ٶ��V= `:w        ���˷�	  S�        �K�KD[�g  LI�        �/}y��  0-�;        �_r�F��z ���         ��� �	�        "����l�3  �&p        Ȍ\_�W  LO�        L���٫g  LO�        �-{�z�^ @�       ����%"�� ��        �V�=r�V�  �/w        `Z��DDV�  �/w        `Jٶ��V= ��        S��K�  �C�        L'�і�  ���        ���v �c�        S�}�hk�  ~B�        L�{; �q	�       �i�~��[�  ~A�        L�{; ��	�       �)�v��{�  ~C�        L �� ���        ^�׈l�3  ��;        0����V�  ��        ���z�� pw        `\���� NC�        ���٫g  �Nw        `L�#�K�
  >@�        ���� �L�        �x�G���  |��        N_^�{; ���       ����yo 8#�;        0���DDV�  ��        �0��ۭz  �$p        ����v �3�        CȾG��� �L�        �߾UO  ���        ��e�"�R= �/�        ����  #�        ���޾V�  ��        ��yo ��        8-��  c�        �� `,w        ��r_�� F�        �R__�'  pgw        �t�� �I�        ���v �1	�       �S�� 0.�;        p*�� �%p        N#��{; ���        �i��{; ���        �)�D��z  $p        N����  x0�;        px��m�� ��	�       ����K�  �@�        Z6��  ��        ����  ��        ��m�� 0�;        pX�� �"p        ��}�� �	�       �C�� 0�;        p8�� �$p        '���	  �        ��m��o�3  ( p        �{; ���        �ad߽� LL�        ��v ��	�       �c�-r�� 03�;        p}}���� @!�;        P/{�v�^ @1�;        P�{;  w        �Z���{;  w        �X_/ѫg  p w        �Nf�v�^ �A�       �2}�D��v  ��       �"�zo �w        �Dn��l�3  8�;        P����  8�;        �t��"�^= ���        O� ���        O��ѷ�  ��        x���TO  ��        ��d�"�Z= ���        O��k�  L�        <Go���z  &p        ��{o ��        ��e�ܮ�+  88�;        �p}�DDV�  ���        �ceFn��  ���        x��]"�W�  ��        �e�� ���        ��-"[�  NB�        <L�� ��       ���}��[�  ND�        <D__�'  p2w        ���m�� ���       ����R= ��        ��=r�V�  ���        �]��Y= ��        w��� �4�;        p7��"�U�  ��        ����R= ��        w��ѷ�  ���        ���  |��        ���{D[�g  prw        ��r}��  � �        ��d��n�+  ��        ���^""�g  0 �;        ��]�G  0�;        �i�-٪g  0�;        �i}}��  �@�        ��d�"�V= ���       �O��R= ���       ����ߪW  0�;        �a}�DDV�  `0w        ��2r�V�  `@w        �Cr["�U�  `@w        �C��Z= �A	�       �w˶E��z  ��        ��z  �        �=r�U�  ``w        �]�v���� ���        ���z��  ���        ��Dd�� ���        �u��  <��        ���"�R� �	�       ���۵z  ��        ���ۥz  ��        �����z  ��        �Խ� �Dw        ৲�m�� �D�        �O�� ���        ?ʌ�n�+  ���        �A��3  ���        �A_/�  ���        �N�-�o�3  ���        �Nn��	  LJ�        �#3r�U�  `Rw        �o��"�W�  `Rw        �o}�VO  `bw         ""��m�� ���        @DD��v  �	�       ��H�;  ��        @�Dd�� ���        @t��  ��        f�[D[�W  ��        f� ���       ��R� �A�       `b��٪g  @D�       `j�]�'  ���        0���R�  �&p       �I�v����  �       ���v��   ��       ����}��  ��       ��r�UO  ��       `B�]�'  ��        0��׈l�3  �w        ���v  �J�        3Ɍܗ�  �Sw        �H��3  ��        0��]�'  �/	�       `�E��z  ���        &��[�  �-�;        L"�k�  �-�;        L ����  �[w        ���v  �@�        �}��   $p      ��*h    IDAT ���Fd��  $p       ���~��   �"p       ���� ���       ��r_#�W�  �w�       ��r�� �y�       `T���R�  �M�        �z��{�  x7�;        *�[�  ��;        �(�w  8�;        ��=�g  ���       `@}�UO  ��       �h�G��z  |��        ��Y=  >L�        ��۵z  |��        F�=�m�+  �S�        0�ܗ���  �)w        �[�  �$p       �Qd
� 85�;        �-n��  �iw        D��	  �%w        BF�k�  ��;         �%"z�  ��;        �-p �s�       ��� �!�       ��r�"�W�  �/�       ���~��   w!p       ���}��   w!p       �˶Fd��  w!p       ��� �H�        pbw  F"p       ���-���+  �n�        pR}�UO  ���       �I�VO  ���       �eF4�;  c�       �	e[""�g  �]	�       ��r_�'  ��	�       ��r_�'  ��	�       �d�m٪g  ��	�       �dr_�'  �C�       �d�  �J�        g�=�o�+  �!�        p"�� ��        ND� ���        p���#  �a�        p�����3  �a�        p�/�  ��        p���	  �Pw        8�̈�U�  ���       �	���g�  x(�;        �@�K�  x8�;        ��ۃ;  �M�        G�=���+  ���        pp�/�  �)�        pp���  �)�        pp�<� 0�;        X�-"{�  x
�;        X��z  <��        ,w�;  ��       �ae�w  &"p       ��ʶGDV�  ���       �A��v  &#p       ��j[�  x*�;        �w  f#p       �ʶEd��  O%p       �#j[�  x:�;        P��z  <��        (=� 0!�;        L�="[�  x:�;        ��v  &%p       ��ɶVO  �w        8���  �I�        G�="[�
  (!p       ��� ���        p ��  �K�        �m��   e�        p���  PF�        �m����  e�        pm�^   ��        p��  �M�        �� ���        � 3���+  ���         ��v  �       �d� ��        �@�  w        8�   p       �z�#�U�  �rw        (�  ��       ���  ��       �Z߫  �!�       ��w  x#p       �J�#�U�  �C�       @��{�  8�;        Tjw  �?�;        ��  ��       @!�;  �C�        ���  �O�        Uz��^�  C�        E�{o ��       @�;  |O�        U��  �M�        E<� ���   ���;�m]ɡ(Z�|���_���C'�-�,i-���`�     PbC�  _�       ��v�cl�g  @+w        ��a�  ��       @��.p ���        P��Q}  �#p       �� �'�;        T�,� �ww        ȶ�?  ���        �mw��  ���        �	� �!�;        $���T�   -	�        �w  xH�        ɶM�  ��        ����  �%�;        d��  �A�        ���G�	  Ж�        2	� �)�;        $���T�   m	�        �f�  ��       @��~�>  ��       @�M�  ��        ��Q}  �%p       �4�w  xA�        I���v  xE�        Y�� �Kw        �r� �+w        H�m�'  @kw        ȲYp �W�        ��.p �W�        �d�>�O  ���        ��.p �W�        �e�W_   �	�        �vcl�W  @kw        H�Yo �]w        � p �]w        � p �]w        Ȱm�  @{w        H�Yp �]w        � p �]w        � p �]w        Ȱm�  @{w        H�Yp �]w        �`�  v	�        �w  �%p       �� `��        2lw  �#p       ��mÂ;  ��       �Ѭ� �[�        p4�;  �E�        ۆ�  �!p       ��Yp ���       �pw  x��        ��o ���       �p
w  x��        'p �w�       �h��  �!p          ��;           -�       �h�V}  LA�          @w           Z�       ����U�   S�          Ђ�          ��           � p          ��;           -�          hA�          @w        8X��>  � p          ��;           -�          hA�        G���   � p          ��;           -�          hA�          @w           Z�          Ђ�          ��        p��>   � p       ���� �-w           Z�       ��L� �;�        p8�;  �C�          @w        8�w  x��        �p �w�          hA�          @w        8ZD�  0�;           -�          hA�        ��'  ��        p�� �;�           � p          ��;        .�  �)�       �h�v  x��        �p �w�        �T  ��5       @#�  �K�        )�  �G�          @w        �� `��        R� `��        2Xp �]w           Z�       @
�  �G�        	"�  �G�          @w        �`�  v	�        ��  ��          hA�        B�  {��          hA�        "�/  ���        � ��  ��        �w  �%p       �w  �%p       �w  �#p       �� `��        R� `��        2Xp �]w        H� `��        2Xp �]w        H!p �=w        �`�  v	�        ��  ^�       @+�  ��        �� ��;        d	�  ���        Y;  �"p       �4w  xE�        I;  �$p       �,w  xI�        i�  ���        ��\  ^�c       �,a�  ^�       @���  /�1       @�  ���        ���  ^�       @�;  �$p       �4w  xE�        Y,� �Kw        H!� �W��        �w  xE�        Y"��  ��       @�� �3w        H%p �g�        �)$;  ���2        d� �S~�        �("�O  ���        �ɂ;  <�        �,� �Sw        �d�  ��[       �D!p ����        UT   m	�        �w  x�o        2�w  xF�        ��  ��        EHv  ��e        �d�  ��       @���  ��       @���  �#~�        �M�  �)       @���  �%�;        $�  �2        d� �C~�        �M�  �)       @���  �%�;        $�  �2        d� �C~�        �M�  �)       @���  �%�;        $�  �2        d�e�a�  ��       @�� �ww        ��  ��/        *� ��d        (w  ��/        *� ��d        � p ���       �@� ��d        � p ���       ��"� ����       ��w  ��/        
��  ~�K       �
��1��
  hE�        U�� �~�        PE�  _�!       @�;  |�        EB�  _�!       @�E�  ��        �Xp �/��       �H� �?d        �"p �/��       ���  ��C       �"���'  @+w        �Q}  �"p       �21FXq ���        P)$<  ��1        T� ����       �P,k�	  І�        *Yp ��       @�� ����       ��"� ����       �R��  @w        (!� ����       ��"� ����       �T�a�  �w        �k�  Ђ�        �Yp �1��        ��"� �1�        P/��  ��;        �E�  c�       �^�x  `�;        �� �C�        �bY�O  ��        P-�1FT_  ��        Ёw  �       @!�  �b        h ;  �       ��E�  w        h B�  ~�        Ёw  �       @� @�        �w  �       @��1��
  (%p       �.B� ���       @�Z}  ��       @!p ���        �E� �6�;        4a� ���       @� �8�;        t��y  �6?b        h"�  \��        ڈ1B� �u	�       �+�  \��        	�  \��        :�� ��	�       ��� paw        �$$=  \��0        tb� ��       @#w  �K�        �D��  ��O        ��� �E	�       ��Xn�'  @	�;        t�Xp ���        �L� �(�;        tw  �I�        �Xp ��        �Ͳ�1��
  H'p       ��B� ���       @G˭�  H'p       ��bY�O  �tw        �H� �	�       �!�  \��        :
�;  �#p       ��b�U�   ��        �Q�!� �Z��       ��X�/  �Tw        h*�[�	  �J�        ]-� ��;        4e� ���       @W� ��;        4w  .F�        ]���  �"�~       ���� �u�       ��Xn�'  @�;        t�Xp �:�        Иw  �D�        �Yp �B�        Иw  �D�        �E�2  ���        ��� �E�       ��X��   ��        ��� �E�       �9�  \��        ��� �E�       �����>  'p       ��b�e�>  'p       �	�r�>  'p       �Xp ��        0�  \��        f p ��        0�X��  �pw        �A,�  N̏        f�ܪ/  �C	�       `!p ���        0�e��   %p       �IXp ���        0	�;  g'p       �Y,��  pf~�        0�e��   #p       ���z�>  #p       ��,w  �K�        	�;  '&p       ��� 83�;        �dY�� ����       ��,k�  p�;        L&�[�	  p�;        �f� pNw        �L,�O  �C�       `2���'  �!�        0�e�  ��/        f�ު/  �_'p       �	�"p �|�        0�e��   ~��        &��  ��	�       `B�ܪO  �_'p       ��2F��W  ���       ���� p2w        �T��O  �_%p       �I�w  NF�        �Z�  ���        &�:ƈ�3  ���       `Z1�b� ���       ��b� pw        ��w  ND�        ��O�	  �k�        0�X-� pw        �Y,�  N��        f����   ~��        &�� �s�       ��b�U�   �B�        �[�  ���        &���. `~~�        pV� 8�;        ���;  �M�        '��  ��&p       �3�� �	�       �b��1��  ���       �;  ��    ����Ǯ��������)�EY6eS�eE�D�X��4
6.p�"�Vۥ��v*��VR��O��-�,���z-k%Q�1��P$[�g�9�{^�V?�H�{9��\   ��w  X.�;        4"��z  <�;        ��w  N�        �p� ���      ��Ml    IDAT @+2#:W� X.�;        4�w  �L�        -�]p `��        А�]p `��        А��  ,��        Z�!r `��        И��	  p*w        hL�� �B	�       �5�� �e�       @c�""�g  ��	�       �9��#  ���        Р���	  pbw        h�� �%�       @���z  ���        ��Y=  ND�        Mʈ~�  '"p       �Fe7TO  ��       @���TO  ��       @���'  ���       �U]�}�
  86�;        4�w  �D�        -� � w        hXvw  �C�        K� X�;        �,3�w  B�        ��~��   �"p       ��e���   �"p       ���c�  8�;        4.�!�B  ,�W�        ��P�   �J�        +���z  <��        V ��z  <��        V@� ��       `���D�  ̛�        V�w  �N�        +!p `��        �w  fN�        +����!  �˫U        X��7�  ��        �&�X�   K�        +�;  s&p       ��~����  �$p       �UɈ~�  �$p       ��I�;  3%p       ���~S=  I�        +�;  s%p       ���.�� 0?w        X!W� �#�;        �P���	  �w        X��  ̏�        �(���W  �7�       `�\q `n�        �R�� ��;        ��� ���       �Zu}D��+  �kw        X1W� ��;        �X�c�  ���        �lp� ���       ��e7Dd_=  "B�        ���X=  "B�        ��öz  D��        p� ���       ��e7Dd_=  �        @D���	   p        "r� PO�        �� �,�       ����Ⱦz  +'p        """W� �%p        """{�;  ��        @D� �'p        ����W�  `��        ��r�VO  `��        �ײ�TO  `��        ��r� PG�        �^v�X� ���        ���;  U�        �7d���  �J	�       �o�a���� �
	�       �oɈ~� �
	�       ���a[= ��        ߑ��z  +$p        �#�1"�E  \,�@       �Gr� ��&p        )�m�  VF�        <��  \4�;        �h]�}�
  VD�        <V��	  ���        x,�;  I�        <V�����  ���        x�̈~S� ���        O��� ��!p        �(�m�  VB�        <QvCD��3  X�;        �T�� p�        �S尩�  �
�       ���~Y= ��	�       ��ˌ���  4N�        K��	  4N�        K���	  4N�        K�cD��3  h��        8�\q ���       �c�a[= ��	�       �c�~Y= �F	�       ��ˌ�7�+  h��        8��  ��;        p"ݰW= �F	�       �����n�^ @��        ��尭�  @��        ��	� 8w        �Ĳ#R~ ���
����       �!#�M�@+@c� 4%#��       k�öz)p�)w �2M�m       E�s��J �6 ڒ�m       &��~S�V�w �"�1�g      �r��i% h� m�:�6      �$p�Z��1l 4eJ�      .RvCD7Vπ��t� �Ń��t�m       �w(��� �,� h��Wo       X�;ԙb��)l ���n      \��ǈt��h% h� mI�6      �
��C� h� ��l      (��^�X��.�7 �YД�&�6      �9�!G�Z	 ��@S��<�       Jd䰩듓� 4E@[�i��       �V9�UO���B+@S� �%c[=      `�����4\�̱z �%�; ��      T�.��T�����x�CW�h������      �BݸW=V�ͧ��; ��      �Pۈ���*w�P/@3� ��w      �J�E�c�
X�m�� �w Z��       źa�z�ʃ]�K@3� 4dʈp       �X�Z[�HC�q��f�h�[��cDd�      ���.����E9�����f�hƯ���7k       3����E針�p 4C�@3��]�      ��nث� ��;4 4C�@3�m'�F      ��������
]i& h���f���       s��+�p:� �Ќ�G.�      �I~�a�e�w ��1�Wo       ���"��z��A�  8+w ���]��       �7�W=��;�; ��Ў�	�      f��p�v�� �w ڱs�      `v�>��W@�v]�; ��Ў��       3��+�p�r7	�h���f�ެ      �P7��\e�WO ��"p�.�      �S�G���ЬGh������      `�\q�s�[�h���v��      0[9
�Ἰ�@K� �ç�      �+��~S��4E�Wo ��"p��L�      f�\q��0M��� 4C�@;��      �X�{��3�Ew �!p�%w      �9�.��T���dN�� ��hF
�      f���'@�:�h�������       <Y{��3�)S�a� 8+w 2=W�       ��Ȍ��+�)��]��  gE�@K�       ��^�hKƥ��W# ��; -�R=       ���a��%8C��_��a� 8^%Є[��W���      �qd���;���W�Vo �� p�	��x�z       Ǘ�����=�V� ΂��&L)p      X��7�WπfS�� �	w �0��I      X���'@3�~�� �	w �0M�M      ���W=�1ew�z ��; M�B�      �4��X=���j' h���&tޤ      ,�+�p6�]\��  gA�@��w      �%����	І����; ��	�      �(��~[��o
� M�Ј��       ��+��즌�� �,�h��      `�r�~y�8�)���  g��B ����^�      ����a�z,ZNӵ� p� ��w      �E�Q��$��� �,�h��       K��&"���\S
�h���F��      �t9�WO�Ś2� 4A�����˥��       �	���2�͍�?<�� �J����_\q�      �]�o�W�bݿ�ߨ�  �J�����\��       ��p�No�$p`�� ,^�\p      hD{!k��麝����J���<r�      ����z,Үs$����x����      �!9TO�E�v;GX<�; ��w      ��d?Ftc�X�k� �Y	�h���       8[9�UO����X<�; ؽ\�       ��Ս���3`Yv�#� ,������	       ���"�m�
X��� �Y	�X�.nVO       ���xP=�e�]��  �J���M�;      @�r�Dd_=�w �O���]�����w       p>rܯ� ˑ�SV� �g!p`�r|p�z       ���I�7?��׫G ����l�N�      в����+`1v��[� �Y�X�)�       ��6���q=|8h) X4�; K�M      @�r�Fd_=!� ,����˗�       p�2rt��c7MZ
 M���yS      �
���%�x�z <�; K'p      X�����W��ej) X6�; ����To       �b�+��T��; �&p`��W/       �b䰍Ⱦz��4ݬ�  �B��b���݋��w       pqrsP=f-C���	�X��>��{��;       �8ݸ~TO��B���P= NK��b�}���       \��"�m�
�����U= NK��b�v��      `�r<�� �6<��Wo ����XSī�       �x9l"��z��ԇ�� ,����ʈW�7       P�s�kw �K��rM��      �J���'x�)oUO ���
���x�z       E2��܁��I��b	�X��w      ��ƃ�	0K��^��  �%p`��|��6"nT�       �P�G{�+`v2��� �� ,�?歈��       �JW�Ủ��Xw )��]�      �z9l"��z�Kƕ�����3 �4� ,�Qt�Uo       `��+��mG�� ,������	       ""r܋H)��.�� �4��`�2�v�       �"#GW��M�
 J��R��      �׺q?"�z�G���' �i�X���       ������+`6r�� ,���Ź��Gۈx�z       󒛃�	0��j� 8�; �����      ��d�����0SN�To ���8]���	       �T�;DDDF܌���O| �8w �{�z       ��^D��3`��n��j� 8)�; ����]�      ����q�z��Ç�~X� NJ����"]p      ౺�ADd�(�������89�7_       <^v��^�
(7��� pRw '#^��       ����z���� pRw �ֿ���)�Z�       �-�1��g@�I��	�X����7�7       ���R��5�nWO ����(�._��       �2��}�(�7�|�Ѷz ����eI�;       ��;+��c��U� ����(ݴ�      pl9�G�L���ؾQ� N�+7 e�\p      �2#ǃ�Pf�t��E��,w�'       �,�� �R�U�$p`Q�j`1��ٯ^����;       X��"ǽ�Pb��� pw #��Wo       `��ͥ���p�r��7 �I�X�.�7�7       �P]9���M߯^  '!p`9��S=      �����	p�2^����J� 8.�; �1E�Y�      ���n���3��僣7�7 �q	�X��V       `ٺ�+��Q?��z ���E�����U�       `�r�Dtc��P9�~R� �K��"|~���W�       `�\qg}��� p\w !NoVo       �9n#ҍ5�#c�S� �K��"Lw       �HFn�G���"o���; �8� ,BF��z       ��ƃ��O����A��z �Wh ,�.�      p�2#GW�Y�i�{�z ������+�^��      @[��ADd��(?�  �!p`���x�G���      @c����W������ �8� �^��f�       ��m.UO�1M��� �8� �^F��z       ����a�z����a� 8�; �7e�U�      �v�+���ҵ�W�U� ���0S�]=      �ve?F���p�2�}G�=�; �v烏��O�w       жn{X=���92��	�����oF�X�      ��}y�}S=�U��� ̞��Y�.��z       ���;����O�7 ������Wc      p1�߸�N���� �i� ���;       �۸�N�2�����+�; �I� �[
�      �89��N˦n�oW� �'�0[7�э��Y�      �u�6��'�9z��  �&p`��ީ�       ��䰍���p.��V� �D��lMS��0       %��+�4j��TO �'�0_]�]=      �u�a�w�4���� �$w �k7�S=      ���6��Ӟ��u���V� ���0Kw>�hoU�       `�r܋��p�r�?rt���0K?�y;"6�;       X7W�i�.�Wo ���0K�����       ��+�4'��w fK��,M9	�      �W�i��v� x�; �4E
�      ���"���gg�~�~�Y�`~��WcF��0       3��m�G���8��o�N� x�; �s�ߊ���       �W�iδ��� �Q� �Ov�VO       �o��6��G���M�;� �Q� �N�$p      `vr��;��Q� x�; 3$p      `�2rsP=�H�U�  E��������       �R7D���˜^������� �m^i0+/u�y3".U�       �Gʌ���6M�q;�[= �M����v�UO       �'�6�Wπg6u��z |�P=  ��.�_e�fo;�q�7����f�c3�1�]�]F�_�	:���h7��n���ރ�q��Q|�Ńxp�+�       ˖�mc��慎�3�I�������|/b����}W6q�`�����	��w1�}l#"�_��{���/��>��~q?&�      ��q/�ާ�Q�8�)�w�7 ��9��l���=�̏#���]f\���.�ǥ�1�^�<<��ǟ݋�|�E|q����"      @��w]qg鎆�ϟ�����g�C �+.�0}���n7��Wn����A\;��R���.�_ُ�W��ӻ�>����޹��      ���q����cZ,V��ßE��� _�0G��=_-�^_��/\ދ����p�?���w�?������c�;      ���0vw?���v���C�����������}/^=��W�#g�3�^�׿x��7���{�-       ���^D7F�TO���x�z �!�; 3�?�^�źvy/n=)�����H���x�ֵ��O�Ư�Y��I      �}y����3�Tr�ީ�  h&wRX���������;�{�!^�q9������������I|z��      ໎>�ǈ���3�4���ϟ�����g�C  "b��RX�a߫���ˌx��A��ʵE������|5n�p�#�      ��t���	pZ�.V= �"p`.~^=��5]ܹu5^~�Ң���ǝ[Wc��      ~/�MD����r��6 �e 31�I��ϕ�����>VO9�1�x�Z���      �F��\=N'���	 ��; ��|��6"|�U�^~�R�v���^v}?�y5���W=      �������Y���w�7 �W�*� X�O.���7�ˌ�/����    IDAT]��TO97��޸/?�z
      0���Ch�޸�'���{��5�����u��޽}������1v������461c443ʌG�0�W#ED��`��H�m����m"�r��͈DJ�&b2�}�Z�V�����E�>�aw�CU=���Hv�v��W�vתU���� ,w @�X�NW����_���S�ų7�+ۑR�      �6W�YJ)�e��S�3  ������WȰߍ|���wk���+��=���      �۵ౕ��ӵ  ����J�� ���A/~�����K��[#w       RӍ�ݨ��%E�p� �0p���_��("������n��^���z����5��^5r     �u�[��,�Rʇj7 @��; �u���j7��v7���.D�xs&"��A�te�v      PQj��z���<R������� � ԕ���������>�b��]����l��       *j����\:��3� ����J����������u��!�{f3.�kg       �4W�Y*%�Gj7 ��; ռ���\����������{����F�v      PI3�3-�E)�'j7 �WN T3o��"<�m)������EJ���nz��)      @���߬]�$E�h�|�[���f�@5%��x|�n�����v��xT�&����      �����"��X,������� `�Y�PM*�˦Ӥ���/D��%���;�ޫ;�3      �R:��(��� �7�4 ������b����<��^݉��'�=�[��za�v      PA�o���RhJ��� �7w �z�߹/�/oǅ�A팥�¥���jg       �.E3��g_N�õ Xo� TQJ��xt]?5)E|�s���x      �&����X,��K������ `}YVPG)/�N��z�x�UWNS��ċ��kg       ���2h:���� ��2p��=s�;"ŏ����5)��>��&�NY9�l��֠v      p�R���B[.�3� X_� ��~���N���KW�c�߭���^�����c      �n��'>��J���	 �/�* �]i��xw�w7��ΰv�J�v�x�7�      `ݤN/Rw�v<TJ�W>�͝� �'w �_I/�N����x��V팵pqk�<~      ����T;�^�n�~�v ����s�̵�\�(�y��Ӥx�s��4�H9//^ގ&��      �JӉ�sŝŕ">^���d����G�������^����?E��m�y�     `�_q7�ba}�v  �ɫ# �W�O�N��v7�qygX;c-]�݈a�[;      8O��4p���Oĵk.�p 8W9��vo�Ӥx��N팵�R�K�������j�   �NJ>�m9�M��"JDD��˓z�Ž��;K���a|�?x�_o�����SDJ��ٻ�����1   N�ߌv:�(m�x��s�����[���b����|��/�(����{��v���R��F/.l���v
  �
*�������˽?%Gyӯ���C�gX|ʚ�C�tw�D�;�O�� ��?����E���  �4�hۑ'�k��[���υ�; ����s�D��ka�iw��v��3��.mŝ���C�   <T���������w�~o��hW�W[����*��}��ߖ���?�0|词�  �I�mDL�yV;ޠI�g#��jw �^�87)�_���[u�ﹲS;��^'.�n�����)   �<0\�m��F����s����������:�O�����9�u��:��1|��b<  ��i�;��7jg��R>QRDr��sc��9))����+;�뺢�H���7_�D��?   ������<^�w}�}���Si���}�O�[��m"��������t\�  VV��#u�Q��)pOJq��+���^�7��n`}�p.�{��~��x�vo��ыg��3x�n��+6�?��N  x'����x�>�7jwy�ww�J��!�[G��d��=�7wG���  �PlG��;<�ݼ�OD�p~�8'��x��"^��];���za3��Lb�~   ��ܿ�o��윏r��Z۾�>=p���|:�-  ��JM7Ro#��1,G��g"��jw �>�89�/�T��]�݈�����Ӥ�za#��Q�  `������!�Kr,��O�����0���{��1��;  P_3؎v6	OAcQ��()"yC�saj��{�z��g�ݏ���)�v������K�E�s���7\q  �^)'����e�y�v�;k���{7R�d����   �)OGQ�^���4i������jw ��m��]�z�#aܾP^��eܾ�&���a���?  ����;d���}Cv��D���\~O���7���vN����  �hz��NǾgga�����0p�\�p�Rz�v�m�qigX;�Gtew#�nF�=�  xL%_co�Ǻ�����x|��CN~u"E�&R�w����<  ��H)��N�ɭ�%%��F�S����V �\*�CV��=W�k'���&.��ۇ�S  �E��7��K;s��E�(m�y{�W'����7�߽I  <��F���v
D��hDI�� ΜwR8SW�}����߆�9���0�{u�v�i:�����(�&   "�/���(�ɐ=�"J�]��to螚�� ���m  <\ig����3 ""�4�������w�; X}.�p�>���I)�{f�vO��m��� n�N  �[�Q��ɐ�evXn%"ώ��<��y`���Gj�F�  �=�Ӌ�݈2��g꛷�OG��; g���3դx����pyw�nS;�'t�¦�;  ����'��{�فՖ���ߟG�{��=p����ݐ  ���w�=8�Op�����"⿮����n( g��_w�M{ߍ�K�S�]�R|�{.E�c������q  �����v�������N��w�яH�� �u���Ljg�������K�^��.`�����y6�$���Ջ��+��;  ,���٧'���xT%�����:�:w/��]y ������F��v
k-�\�h?���.`��pfJ�WRy�g�Ӥ���Q;�Spqk�ib޺�  ˠ��7�� 8M��2o#擓���W����wW� `u��`;��v��\��Sa��3p��4�|ƾ���6]o_)E<�=��n�N  ޢDi��>�(>�
��������ԉ���Gө�  <��ۈ��#��>SO)�r� V�gUp&����Ws��aY]Q����}��4�䯊ɴ�����Q;  ���F�O#�YD�.u"u�'�� `�vy�_;�5VJ�E�u�ƿ�Wwj� ��\p�L��J��ڞ��iܾb��Nlo����U  8w�=���,��F�F��<.u���w�  �$�_���'�SXS)�^�g~."���- �.w �Fi>QjW��n���;������Cw  8%�#ڙA;��Je���4�{��S��ܯ  �E�v�����SMI�w ΐ�; ��G��u����t�uwyw���+��� �v� r�  ���O.�_i���.8_y%ϣ��ǿnzo���  ��D�oE��.am��k �ڜ� �Խּ�rD���Xg)E\�٨���4)v7��3  `%�v�� ��h�����Ӹ "Ϣ�ƑoF{��h�7"OGQZO� �ښ�VD���`m������׮ `u����K�sW��K;����*{fg�FG�3  `����J�Q�vQr�"�%Q"����C#"R�ӿݽ1� �s�R4Ýȇ�j���J�s�LD�O�K XM� ��R�/�nXwWv]o_u;��v����8  �nJ;;�Ϗ"��� ���(�I����שs<v�#u{��� �:H�aD��Nk���R*�w Έ�; ��k��?+�W�c�]�İ�b֪K)bw�7^��N ��S��+��#W��Ci���Qf�h"u]w ���w#��#�s�9_%�/D������kj �bR�s��������[��	  �0J;�<E;���w#ފ2;4n����{�܎v�Z����GQZO�  �Ӗ�n���SC�z��� �&�8U%�����A7��������~t�m��x  �Q��Σ�O����� x�<�2�E�D����{w�ۏ�T�  �^3؎v>�A�]��~)"�m� V�� �����g#�õ;�����8G)E�� �:)\~�����(��q;�2)9��0���㿗{�  <��D�߮]�z�D�  V��; �&���זj��&.;����~�  8[�=Bފ���!dB,�>�t��h�7�L���  �R3��o�[��g>��/Ԯ `�tk �:R�_�H�z��D�?�����GJ��. ��S�<�le~�g�s 8/�4r;�8���"�����H�g ��h�;��7jg�FRJ�No���k� �Z\��T����lF�O��Xg�v6j'PA�I�5t� ��W�<��A���ȣ�(��v�u�gQ�^�<�;~���N��4"|�  &u���~n������ ��q��S1ߜ&Jڪݱ�����;�3�dws��?  ,��΢�'Qf�����`Q�6�le6�H����a�n�v  ,�f���("r��D)铵 X=.�p:J�B�uvigX;��v6�0 ��Q�i�ɝ�k���(ӑq; ��d�oܿ����?  ��t"ܦ���T�s����Gjw �Z\p��}�;�t��E��Ӥ��5��AE�~'z�&f�+  ,��N��&Q�G�� ��7_v��/�wz��  ������0"�k��&J�."�}� V�� <�go�/���XW���4�v�mm��-  ���y䣃�K�7�Ǉ�� ���F��"��]v �H�vkG�FRI��n `��p
�j��K;��	,��~�  �?j�E�E��p�N.���~����GQ\� `ͤn?R�ϒ9'M|����/�� `u��t�_o"�/��XW�nl��3X �C� ��mG�F� ,�<�2=�<�;�OG%׮ �s�v�<��"�ݍ���; X^� �T������jw���[��	,�A����v  ���#OG�CA�v �E�E9z=ڃ�F;�evh� �jk:�[�+X95� �+( �Jj�j7���<`�w  �T�2�D>���kQ�^�ȳ�Q �d�i���h^�|x+�|�v  �����x*8g/����8�� �>_;`]m�1�ujg�@6�  ��2? �n �*z����N���  X%)��n��AJW��L|�v ���� xbW�}�Ǣ����XW]o�M\p ഔvevx<f/�v ������Qf㈦Mo#Ro�܋ `��n?Rwxr� �N��+��� `�yG�'֤����w�d�ߍ&��  ,���L�ю�#����}�� ��<�|t����'�  ���n��q�R�O�n `5x��+)~�vú�tc����`��t��  <�e~������ND�Վ�R��''_+�"O�D���Q  ��Ri�U��U��/~���jg ���x"W^���%~�vǺ��z;a� ��(�,���Uڛ����(m��8�h/��(�CO; `�4�͈��9S���/׎ `���D:���nXg�y�a�R  <Dɑ��hG{���Qfc�< xR�4���ɇ�nGi���  ��h���#Xq%���n `���DJI�V�a]���:�3XP�  �I�O#ފ��(G�G�y�$ X!%��0����Ȧ#  `��N?Ro�v+,E|��Ǿ�S���f��c�������jg�W;����FJ�+  �.����^�|x#�|�v ��<�r�����[Q殺 ����ND2㌤ƅ�/�� `�y��ckr�V�a��l�k'��R��\q XO%�|��f���k� k��kr><��^���f  ,����᬴�_�� �r3p�	�/�.XWMJ�5p��w6�uj'  p�J�G�ܹw-6ڣ�I �]y������N�<�]  �z��8��OǇ�n� �3p�<��~2"~�vǺ���iR�ܠo� ���(���ȣ�(�qDɵ� ���Qf�ȣ�hG�Qf��;  u5�݈��gN_��x�ʳ�P���e��cɑ��nXg;�>Aϻ���  8+%G��N���t� �Q�E��v� ��RӍ�߬���J�/�N `y��J��mox��n�s� `Ք�4��h�������N �Vy���f��� p���vD��E��gk ���xdW����"�}�;�U���F�en���� `5�e:>��~#�|R� 8+�Q�Û�_�����k �.R�f�S���Ry��O_�p� ���; �,5�˵���f�vK�iRt;^� ,���"O�D{���k� �NJ������;��   �^�#u��3XA%ů�n `9Y>�h^�ލ_���ζ���	,�^��< ��RJ��a������(�qD��
 �+G������V���v  +��)�-E��� XN^� �H�\}���l�u�9��N`�����	  <���'��_�<��g�� �S�ȇ7�߈2�DD�� �*j:�[�+X5)����W�v ����G�4����Ӥ��yt}� X�2�D;�y��Z; �h�i�ɭh�"OG��  NW�ߌh<Y�ӕ�ޫ� X>�O ��?���(�˵;��Ơ)ծ`��\p X<�D���Gi�[�v ��J�����w��y�"  VF�f�[;��">_���c���j���#b�v�:���<����2 `Q�<�<���k���D��v �r��8�h/���(��A  ����E�m��`�4��~����� `�X>��R|�vº�tk'�dz�  Օ�4��ȣ�(�qD��I ��j�"ތv�e6�] ��k;��95�i�# X.�O ���\�.��O��Xw.��:�T; `M�(��hG��oD�� �(�"OnE{�Z��8"J�"  �QJ�wkW�B�H��� �r1p�Mc�jD�kw��^��^חl��  ����Q�{�'�#�v ��J����k����b� ��I�A��v�"�O<���S;��a��;K��j'��-��y�N�w �3W�<����ԣ�#J[;	 ��F�D{����=�. `�4�݈d^�i(Mt�֮ `yx�C]��_�`D�H�u7�wk'��w �3S��ȇ�"������** �����}/��ND��<  Aj��o׮`E�h�P���a���u�W#�B�����;O�i�� �T�ev�h/��(�I�" �ǔ���ǯg&���y�   \�oFt��3X)Ň/���T���`��C��J�r�
\p��u/�  NEɑ�^���ȓ��` ��;��^�E>���� `�5��p�S�)�ޫ�# XVO ����/_���ݱ&�]_�y2M�& ��(yyr;ڃעLG�k' ��2�D�G;����� `����U;�U���k' �,� x[9�Wk71�wj'��:��; ��(�,��ȣ�(�È(��  �^{y|#��Cw  ޢlE4�>��I)>z������3p�-���?ۊ�_��A�F�<9� Ͻa�x?�|R; ��vj� ��H�/Ԏ`�uJ��v �����(��_����D�y
�� ����Q����  2t �MR���Y;�%�D��j7 ���x;_��1w��y; �;)Qf�ю�"ތ0� x{��  <��D�N��Y*?y���3 Xl� ���k�~)Ry�v)El��4,� ު�(�q�{�'�#�v �r�7t���ծ ����^�]�rKm���� ,6w ޠ��W#�ǭ��׍d��SH� ����Gю^�|t'����  �S{y�o� ��R���Q;�eV�k' ���x@I%�wjWplc�z;O��R; ���F�܉�`/�� ���E  ��� `�5Ý�dzƓI)~��O��kw ���� �.��]    IDAT���>�������;Oɾ Xc%Ϗ��(�qD� ����{>�e� �NR�`�vK�i�_�� ��2p������nྭ��;OǾ XG%�#ފ|o��U �y(�����vDnk�  pRo�;������� ,.w ""�k߹�Z��c)E{�<�R�� ��q|����}>�� ����0��^�ɝ��):  ���F$4�@���?�P� �W DDD/�#b�v��n4M�����o �Aig\l?�� @DD�(�q�{���Q ��R�`�vK*w���n `1�)�߭��}��yz%�� X]%Ϗ���}� V�2=�v�Z��(��U  +)�6":��,�r-�# o� ����GK��>-����;O�a, `��b�a; �r(9�����E�y ����N���R�K�?=��� ,�* ���?���m�yz� �*q� `�6��V�#��  VMj��[�3XF����	 ,w�5��W�|PJ���ܗRİg���+� ��{�v� VG>~*O;���ծ ��4���N�v��W����d�v ���`ͽ���Ո�R����n4M��  U� ���(�x?��(y^� �S�^�4K�����jg �X�� Xs����n��6��s:rv� X>��� ��2�D�G�܉(�v  O��Dlծ`����f� ��;��r�/(��x��h���Sb� ,�{�����  k�D����E��"�{[  ˪�oEt��3X*���}����+ X� k�I��""����6��	���� X���.� Qr��ף��# �2�/�i�*�ԛu�/�� `qx����ʟ"�Wjw�FMJ��w���WJD.� ��m���v  ���!��(y^� ���t"�jW�DR�ߨ� ��0pXSwv��"�j��hs؍�>��͹v ��+9��A���(�q�  ];�<ڋ<�Q�� �L��VD�_;����+���Վ `1���߫�[mz�X��v `����E�D�,  <�2;�v�y:
�% �G3܍W�x$���# X� k�W�����X��jsЭ���p� X�D���/�O"��  �P�Q�^�v�e>�] �#HM7�`�vK���R�u�F ��Q.���H/$�9-�	w ��r��f9z=�� pJ�<��h�7��y�  �E�ߊ��kg�R��.z��; ���`ͼ���_���[�{��u}i�t�� @Eev��^������ `U��ȣ�ȓ;>P	 ����n��ǣI�S� ���� ��Q^-����6��	��\���W�Gю�� 8We6>~r�t\; ��HM7��N��AJ�|�c����3pX7)�~����W;��; p�J;�v|#��͈<�� �:*9�ѝhG�QZ�I Q�oFt�3Xt)�۝��kg P��;�y�7��R�O����m]p����G2 g��y��[����v  D�Y��ݧ
y� `�t6.D$�5�Y��[� �˫�5RJ����&������� g�ް}�e>��  oQf�ю���k�  ��D3ة]��K)}��g��C�; ���`M<�ϯF�k�;x{[�^�T��U2�� g���G�G���  ,��#OnG;ڏ��j�  p"�6"u��3Xl���ߩ@=� k�D���;��5t���5�� �i*�/`N"�� �G�g����'�#���  A3܍H�k<\I�7#���`M� ���u�4������9m3��SRf�h���  Xz�>�9;�� @j�G��)��\ze��� �a���M����[����R��[;��fWU��S�Y���'�"J[;  NGɑ'���Gig�k  �Z�#u7jg������� �a��J�o�n��6�h�T;�RJļu] x2%�#ފ<ޏh��s  �l�Y��' T�w"R�v�D������� �?w��«��@�x�v�5��N`�� O��ȓ;�G�Q��5  p.��������  u�&���,�T����Wkg p��V\[�?�����;�mf� <�e:�v�e6��R;  �Wi��btx+"��k  �N��#�6kg��R�|�v ���`�]��?ߍ(_���;3p紹� <�2�D{���ND� ��V��k��q� ���v"R�v�郗>�?];��e��º���#b�v�1�F�q`��e� ���΢߈<�Q\� ��r�;юoD���1  �#�h6.֮`A����n �|���k݉H�_;�w�z;ga67p �^��ȇ�"��#�i�  X\�4�h?��AD��5  k!uz��۵3XD)�x�c�ܩ���1pXQϦ��G�������l�k'���殰 oRr䣃ȣ�(�I�  X%�� ��~ 8�`+����Y�iw�_�]��1pXU����	���\p�l�����a���(S�' ���y��ȓ��� �V���B���fMi�V���� �
���_��H�3�;xg��^t�T;�4��! Q�Y�F8  pj�?<�H  g��D3ܩ]��I�᫟������0pXAMi\o_���s�Jq� �^n#ގ<ޏh��k  `��6��ȇ�|� ���F��v&���k7 p>�V�s_����j����F�v+h��(�v PG�|tprQ�v  ��2�D;ڋ2�� �4�݈d��}%�K/~��f� ΞW  +���DĠv�Ӥ�����s� �S�E{�ez�H ��(9��v�㛮� ���D3�X���".N��Wjw p��V����?#������m{�R�
V�t�i �NJ�G;���fD�A7  ��=r� ���n?R��n�K9�^���g��BG�������mo�k'���3�6 X%G�܉<ڏh�j�   '����-�� NY3؉h��3XM�ЕO��O�� �l����כ������lo�j'���sw Xuevxrr�v  ��2��� p�R�fx!"<&�c��|�v g��`E<�7W?�">P��w��4����r��l�: ���N��G��v  �k�  �.uz��[�3X�.�|�b� Ύ�;��(�Ok'�h�\o�Mf��	 �i�m��[��7"�v  ������G�Oj�  ��f�����`���گ�� ��������?�~�v�fwsP;��sq� VJ�2�  �2+'Xu� ���/D$�7"R��k7 pv|�XM4߬���I)b�w��d��N  NIi�юnD>�F0  ��\s 8%M'��n�
A�>p���� �w�%����GJ�gkw�h6��v|��l���+9�����yV�  8Mw��OnG�R� `i��0Ro�v��I��v g��`��N��""�����n�k'�f��	 �S(��hG{Q懵S  �3t�;�� ����nDӭ�Ae��/\��?~�v ���`�]���"�K�;xt;��� ��J;�v�r�1��  �Ci#�oD>:��� [J�/�{��-E�s���� �>w�%�I��D�����u����9g�p�; ,��#O�D�G�Y�  ��2=�vt#J�� ��J�^��v�*kR����jw p����3׾s!"���<��M�OqvJ���]p�eQf�ю���ƵS  ���,��F���  W�ߊ��Y�ZK���̗kg p���T?�߈��;xt����sv�fmO2��W�<��ȓ�%��  F�|t'��-�+  <��ƅ�ԩ�AE)�7j7 p�����_��A����<��"��������G�B+%��A��~D;�]  ,�2�D;ڏ2�} �#KM4C��Z�>t�S���3 8=� K����W#��<��a?�&��`����	 �C��Q���(Ӄ���  �]�6��ȓ;�{ �G���H���T�6�?�� ��1pX6ׯ79�?��������N`�M�`��6���ȇ7#���  ��)�q��Q��7 <�f��x���ʿr�S��� �w�%���\�|��@�υ�A�V�x2��  �S"D;ڋh�j�   �,�"���LǵK  �@�f�B�ĭ��R/���� �t�j�lJ���	<��A/�]_r9;9���]��EP�����AD��9  �J(���D>�Qr� ������%w�Sʿ󾗯kg ���� �ȕk���ӵ;x<�]o�lMf�(�s PW9�ڞ��ٓU  ��W�hG�QZ�s  ���ۈ�ݨ�A)]����v� ���;���g�x|����	���Ѽv ��2?�v�wr�  ��6��F�#�  ��f��tkgPA�� xz� K�W������<�a��^�v+��� �(9��v�Û��]  ��ez��fDɵc  SJ�l\��T�����+����kG �t��D��'�;��sqkP;�5p85p��Vf��W�g��S  �u�E;ڏ2��. XH��F3ة�AmJ��v O��`	���>�J\��������N`ŕq4u1 �K��h�7"On��  �W�ȇ7"�. XH���;���9kJ�������� <9w�%�F�������ub�߭������K�� k�D��"��#Z� ��R�юo� . ��h���S;���D���3 xrƒ ��o�?J�z��ŭA����Ѽv ���΢݈r�zD�`  ���i���(s� x��D�q1"R��U�ڋ���Y��'c���R��ED8��.�s�� pfJ�|ty��g�k   �]ɑoD��	� �/uz�۵38G)ť�Y��� <w������(��<�^��́�%p�&� p&��������v
  �c+�q��%�N XM+��P�:i"�Q��'c������K��휃R"�w 8U%G>���fDik�   <�v�h?J�T  wu6.D�N��KJ?|�S��� <>w��������߬�����=���8��#���Rf����I�  ��Q������{�=�����|�{fzf�\�93����J\,[ #C�1ج�����肍��H8B�J>��#�Vk�S�8IU*��W�*c�C�r�J*N�S`�d�����t�t��������sfz�ӗ��/xVmU������ݏ<�. ������t	W%��J� ��;��jZ�xDtJw���;�X]vx��w:py	 &��W���)]  0a9���h�GϾ `���R����\�TUo�y�co,���1p�B�=����Kwp>ۮ�sEzg� pQy�j;  ��u�n�f\: ��ji-R�o��!WMt ��`
���C�T����Z_.���p� .��W����  �Gs��!_ ���V6"R�tW ����o���� �?w�)s��O�*"}O��gu�� s�F�&Fcc< 8W� �������ȥc  �IUTݭ�H�K�d)b)uW�f��;��i7�c���r���rz�z; <0W�  ~G����� Xh�Չj�Z��@��}������ �w�)r��<�PD����OJ[k�\�Ӂ�; <W�  ^@=���n�ڿ7 �+-�FjwKgp�ҵN���� �w�)�j��5ͨ����}�r5��>5uԽW�  ^L����G�K�  S�lDT��\�T���ȣwVJw ��� �����s��/���m�����h���t L�<�G}z7�>+�  0�r4��h��K�  \����n�9ݼ˷����-]���0%R�>��Ϭ*��\3p�j��Ƒ�� /��W�G�j;  ��ʣ^Խo� R��Q�\+��e��co�U:��f�0~�S7#���3lcm)ZU*���蝍J' ��r�  ���aԧw#�� X<�Ӎ�q�p�U)}���|G� ^��;����"b�t�w�?p�:'}?,��h�{���  LB���DJ�  \�jy#��������� �4w��n����H�-���-uZ����-W�ir�������a�  �9�D�?���t ��J)��f��ͳ�7�r�[KW ��|V������������	,���8��Kg �t�ύ-\m  �4yxM�0¿K $U��F�̫���n ���t��O>�W���پf��չ�w� ""�x�����A�  ���ǃ�{�M]: �ʤ�r����\�TUo�y�co,��3p(�i�߈�������R,�}�ruN���	 PV������Gd�
  �+ӌ��ݍ<v� X��zDk�t�"WMn�p�
 ^�E@!�����G�w���b���������; �+�ύ)F��)   �)7�����. �2��fDj����T�m۝W�� �K��T��>�gZ�U�ƪ'��:'�a�\� J�ќ݋�w7���  Xp9�ٽhǥC  �F���nED*]����i�_��/eX	P��w=�D��^����^_���W�����v On�Q��Gv  `��Q/��A�� ,���D��Q:�K�"ߵ7=~�t �g�P@�T?�yׯuK'�`N�� ,�fx��݈�w   �T�Ϣ��G4u� �K�:�H;����u���� ������;?�G#�7���b�V:���*����ǥ3 �j4uԽ��g�"�%@  ��֌����p2 0������S:�	K��K;��o�t ������H-���]��R:�s2�� �!��Q�ލ���S   �_���wy|V� ���hu�"���\Iig����� �.ߴ W�ֻ>��#�7���bڭ*�֖Kg�`���� �s�����("��5   <�&��A4g'�C  .WՊje�t�R�y�k� S���ܹS�\�x�.������T:�s�3p`~�� ��g"��S   ��<<�fp�t
 ��I�H��Jg0A)�C�K�{Kw �,w�+����zOD���\LJ���*��F1�]�`���8��aD�]  0/�u�0"� �ZZ�Զ�+U|�w��`�p~�N��z��X]��N�t���v �Pn�Q��#�z�S   ��YԽ���.] pi��͈�S:�	I)>�6�_� w�+�{X����;�������0_��i4�w#�Q�   .S3z����� ��J)��fD2ÛU�?��[*���|�\�G���D�����;����7Wk8nb0�� ���M4���g�"�k�  B���D;� ̧T��Z�*����*�z������ ������z���_Y������-��:N ����aԧw#��S   �rM4���# �)��"-_+����*�h<z�]�`��\���'�#ҏ����ZU�����,�{=W� �u9��q4���\��  ����0����!  ��ZZ�Զ+�)������� Xd� �������\����hU�t�ir��G�3 ��r3��t?�W:  �)��'��Kg  \�je3���`r��bo�U�`Q�\�{O�"��WJw07�uK'�������\: �%��ќ�G4�  ���M�0"��' 0gR�Vw+"��ͺ*�/�q�u�]�`Q�&�$���fD�����u�be�C�\��ްt <��D�?�fpM�   �T��D8� ̛���VDxK����C���a�p	v������77]o��{� ̘<F}z7�xP:  �YP���GdH �%��"-���ࢪ����{O��Ed�pr���3v.�,�ccu�t�w6�Q�G fE���$��~D�K�   0K�ѳK7��%  U-�E�8�7��P� �+�`�n�}�OD�7��`2v�VK'���N]o`6�f��~��I�   fU����G�G�K  &�Zو�:�3��*�ޝ���Jg ,w�I��ǭ*�GKg0�v[k˥3XP��g� �e�� �����   ��M4���c�? �y���݊Hfz���Zq��j�������_���.��d�l�FJ�+XD��QGu� x	9��q4�ÈhJ�   07�h��ǃ�!  �S���nG���J������� ���`Bv��X���Z�&�U��qm�t����v �Wn�Q��G�J%B�8    IDAT�   0�r4��ȣ~� ��I�NT+�3�����n X$� �R|0"*��d���FUyz�2�z^��tʣ~4��ͨt
   s�� s%u����Jgp^)����~�w�+b�07����#��Kw0UJq�Z�t�w6��.� ϗs4��hGє�  `A4��h�NJg  LL�|-R���gV��q���
����V������ؾ����H�8<9+�  ϓ�qԽ��cW�   �zyxb� ̕je3����|��ƛ��*��� .h�=�xC���;���"v6]o���Sw �G��9ݏhF�S   X`yx��t �d���VD2ݛE�����V��y�[����\����r,w�礌��(F�t D�M�(��QD�n  ��<�E�?��\: ��VTݭ�H�Kx@�J_�}�U�_�`��\�λ>��H��L�Ζ��sx�z; ��zu�n�q�t
   <O������ZKQ�l���R���#��Y)�0���k��RN?]:���X]���N��ᩁ; e�a/��~D3.�   /(�Q�#��; 0�R���Z:��Rz��J��� �����n��}_D���Lέm4R��`�qS:�E�s4��hΎ�<   �^}u��� ��ʵ��r�P���;��o�t��2p8���'�s�/����Ni��PJ�GQ�>y<(�   ��� s"E��Q�K�� R�����/�0���#����Jg09��SR��'� \�<�G�ۏ�u�   xpF� ��HUTݭ�d�7SR�?���ǶKg �#߈ ����^�">P���q��Ҏzg1��� ,���8��QD   0��aԽ����X�ٖ���#�H�S�O)���Z�� �����T��X)����Ni�� X �G}�y�+�   �ь��� 3/���Z�(����⽻o�Э� ������{�[#�w��`r\o��q�Ľ��t "�Ϣ��G4��)   0YF� ��H�n����ܷt�^j�t��1p�_��i�?_:��r���N�"�� ̿��I4}?�  0ǌ��9Q-�GjwKgp�r|����<R:`��ܧ��[��_S���q��i�oP:�y���{��'�K   ��� s��nD��Jgp?R��r��� ����>�r����?V���r���zg�ǥ3 �c�F}z7��N  ��c� ̅��VDj��>��}�m�=�; 慁;�}������;��ۙ'��py�M� "ץS   ��� � UQ�n����K)u����; �o>�������F��P��ɺ��V:��s���Y� �Q����9;��\�   �1r �@��Qu�""�N�e���Ν�?��� ����eT)�|Dx���Z[���v��q�,ƵU ��\��>}&��[B    "�����: 0�R{)�������8w\q� w��pk�w�o)���q����w�z; �G�hz�.�   ӥF�?0r fZ�t#uVKg�2������}��Kw �:w��ʽ���U���L֍�n,w䧬q��q���I����E���   ����^r#w `vU+��+�3xi��T�t��3pxô�x����LN�J���if�ۿ7p(���MԽ�ȣ^�   �~�Y�=#w `�U�͈�R�^R���o��;KW �2w�p��O�*"�p�&kgs5:m_}���q�t s ף�O�F���)   0;�h�Ga� ̮��VD�.�K�Z?���$�9Y���v�~."���#�V;���ǽa��M� f\����G�t
   ̜<<7r �Q��������U����|��Jw �*�p _��;��c��L֭�kQU�t�]������8��Ks   py<x��k �ٔ�vT�툰��Z)}x��.�0�����?n59�|�&k�ӊ��+�3 ��&����3 �U���wy�+]   s!����Kg  �[ju��n���E�7[���Kw �"w�/����O"�Jw0Y]_��e����~d�v8�\��>�Q{P
   &)�z�OKg  �[j�DZ�V:�������ï*�0k��s�;�ܭ"�F�&ku��k˥3 r�ؿ7(��ʣ~4���\�N  �����Ezc 0����H��������~�t��1pxN���ۥ;���o��N���8<=�qݔ� `��hG��"�+@   �25gǑǎ�  ��Zو�^)��I�=7���?P:`��D�����]����Z[���N��������	 ̒�D}�y��   �J�?�<��  8����Z*���j5���� �����;�鉈H�S��*��}��v�C8����t 3"�èO�F4�;   �j�h���k� �*E��Q�K��ER��t���S�; f��;��vww�)�P�������r�U:""����p�M� "ץS   `A5��"7��!  瓪hu�#�i�ɹ�h��� ��b�B���'^�>R���괫��\-�Q79O�x99��Q4���ȥc   `������ 3�jE����)���~���-�0|����ߍ���L��7֣�R�����{��CE ^Bn��D�K�    �����)] p.�Չ���S%ŝ���\mx����}�o�H�Q���Z�vbkm�tDDD��;�� `��z��݈zX:   �b�8��ax� 0�R{)����|���+;�?R�`���{�)�t��ҳ��aZ���h� /,�Ͼ�<{�9   L�zM��t ���N7���|�����<�#�Kw L3w`!���㵥;����.�Kg��p���O��F��   `��� ��q� �s���"-����wm�++?^:`����>�U郥;��v��[[��3�w��G�?�� `��M�0�ٽ�%   �ȣ^4���  �V-_������R������[:`Z��j������L���k�n�Zcz�����MԽ���A�   ���=� 3��nD�Lf�A�Xʭ�S�`ZY����o/��du��q}}�t������ްt S$ף�O�F4��)   �4��ȵ���Y���݊h-�!"R��v���?,�0�܁�q���ZN�o��`�^qc=R*]��i���y4������)   ���h���q� ��Iύܫv�"���g��{�8 �"���H+g="^Q���ھ�k+���;F�&O���g5g'�#"�N   &%7��"rS� �|R��vDj�.YxUJ_��ʯ��� ���X��>�5)�Kw0Y�V__+����q?�# 9G�;�<<)]   \�\G��P; 0êVTݭ0!,/��C;����� �ķ� r���dD8�=g��햯2�G��ؿ�z;����8��݈��t
   p��a4���  �Z��V�""�NYh)��fy�'Kw L����n�ňxo�&k�ۉW�X/����� �N�Y����"r]:   �
�8""R{�p �����Վ<�[wQ)�a�˾���ͯ}�t
�4p��k;{O�N9�T�&�J)^y�Z�x��#>w�+�@Ayԏ�w���)   ��Ó�#o� fWj�D��Y:cѵrg��KG Lw`��T},Gl��`�v�Vc��%$L���A��� ��9;�fp�t
   P@38�\�Jg  �[�D��Q:c����[?�]�; ���;0�v���?���t���Ԏݭ���<9G<}�z;�b���"OJ�    E�h��M]: ����j�����I��>�u?`,<w`.���_��|�t��ʛ�R�
x���AG~� X8���wy�/]   L�\G�?|�*
 �����#-���XX)�Wvn=^��4w`.����L�*��d�����J�t<��� �)7�{���t
   0M�Q4���  R-_����XX)������#�; J2p���'�`�齥;��N����{B��sp2�3��J���G4��)   ���A4g'�3  .�Zٌ�^)���R�V���� %����;�&�"�U:��z���hU�t<��� �'����"rS:   �byxy�/� p!Uw3��\:c!�������� ��s���ΏF�ז�`�6V�bs�LL���3��Hsv��+�s�   `4�����t ��hu�"�N�E�r��swl<�����;���W�>\���jU)^q�Z��9G|��t W"G�?�<�jq   �A�h��� ̶����m�^BJo�~��Jg �`�̉�R����n�&����u��q�`A�&��A�W�   ��{�p �LKճ#��*]�p������m�� �j��\�y�'�7R~S�&�Zw)n\[)�/���^� .Yn�Q�ލ���S   �Y֌���  ��TEk�����K����/]p�|� 3���<u3�濍���-LN�J񚇶�U��)�%O���K� �,����"�+�  �	h�)Ej-�. 8�TEj/G�j�R�˯���~���ߗ.�*.�3oT�����;��WܼKm_SL����0��xM߸   ��|v/���t ��������d�qURJ����xD�	,�2�L��{�m)�ݥ;��͵��^_.�/���,�q� .I�����#   �eh�G��� ̶T���n�_���7�x�G��� W�70��SO��*=Q���j��xō����r�����3 �$��8����   �\k�}�>{� �m��yv�n�x�~�ڛ�Q:�*�vfָ��D�xm�&�7ף����tz��Q]:�����#�z�C   �EЌ����  ����D���t�bHi��j��� W�U: �<n����9����\�Z_���k�3��M���q4�� ̗�<��r}V�   X$��c*��T8 �bRՊ��D���*�*�q��������v���d
̜�x�/,�����\鴪xō���>wԋqݔ� `��:��~D=,]   ,�<<�<��  ���^���.�_�VT��wl?���C�9����Z�x}�&�;ע���t����a�t ��QԽ�͸t
   ����qd�> ́�^yn�ΥK���o��� ��#S�L��{�kSJ�kDtJ�09ׯ�īv��΀��gN�;����a4�È�f   `
T�h�ވH~� f_���Θ{9�3æ������.�p��fǣw�)�/�q�\鴫x��z�xQ�a�����E����q;   05�� 07R���F錹�R�\��?]���3cww�F�7��`rR�x��F�*I�^�=8��KW 0	���s?�`   �K����  ����i�Z����?�͏K���`�̄��|����L���j�w�gz��FqxzV:����#OJ�    ��|v/�ؿI �ZZ3r�t�ʭ��bo�U�`�܁���v�_����)L��J'nm��΀���}�r f^�Q�#�z�K    ^V38�h��  a�~R���G_��Kg L��;0�n��~0����;��V��ջ�R�xqǽa��G�3 ���D�?��]>   fDn��F�\� `"�ܯ@��k7����Kg L��;0�n���刏��`�^�s-�ھ��^9��0�ru� ��.   x0�(��q�
 ��1r�\)�ͦ���Kw L�u!0��ܩZ��#b�t
�sc��k˥3�%=s܏�p\:�s��8�ӻ�7q    �)���b 懑��J)��ƛ?��� �b�L���������L��R;��V:^Ҹn���^� �)ףhz��.�   p!��$r�~ `~�_��������! ��* �Bn���_���/#�S��ɨR��<�Km_=L�O���� �(��hz�єN   ��<F��F�T: `"Rk�������S�O���kۣ����_-�pQ.���Ν�ʭ���)L��7ף��.�/�?���~� �!���¸   �+����t	 �ĸ�~yRj��[~�u�; .���:;���_���t����7���΀���'��F 0s��z  �yU�9;-] 0Q��Z�����'�J��'Kg \T�t ����'����X*��dt�U���fT�Wg2�N��sG��̚��$��^�   ��U#�:�*o� �Gj?7��eC�MJ�t_��?���_�?J� ����ɩn�/G��3�DJ��ڈv��ӭir|f��t �9�y��   X��(��Kg  LT��i�Z��Su>����� 8/�C`j����_N�t�����X]�΀���Q/F�t �-G�?�<�jn   `��&��aDΥK  &�ZZ3r�����r��\���j� �����O�6W鿊���-L���r<|�1~��٨��z�^�9 `F������t	   ���MDΑ�˥K  &*��"R����S�GJ_���?�/{�����t
��r�(�Ν*W�#�zN,wZ��O�2>��k7 �!7Q�"��%    ��Q/�_: `⪥��V6Kg̓�T�/�z��J� <(w������#�)��dT)�#�6�U��)�N��8:5��	���w�j   @D4�����t �ĥN��}�R�׌�ʏ�� xPև@Q��>�����ˈX)��d|٭��Z�ZL�_����b0�N��|~����   �wT�h�ވH~� �O�E�7�_T�yT�?��?����t��r�(��;��?
���qs�k�����Qϸ`4uԧw��   �X3�fp\� �R���s��=�wQ)�N^j�b��J� �/w���[��)}}�&cu�__/���lT�gz�3 x�G�ۏ�u�   �����ȣ~� �K�:+Qu��'"�7^?�=?T:�~����y��oLM�_"�S���k����WlG��)f�o|�(����3 x	�E�?��M�   �)WE�v=R�. p)��,��aD��)�-�ɸi�p�O�ߔNx9���������rj���s!��W�^3ngf���L9�v   ��D�?��_ �|J�娺����Xo���� ���r���?_]��ɸ��׺K�3ྌ�&>�Z:�����hz��    �Esv�t ��I�%#�	HU�7������ x9>�+����o�����h�n��6V��5�7Kg�}�wO���Y� ^��K   \L����R: ���zM�0"K:�����W��GJ� �܁+��zj5���q�\X��ջ�3����� S,���    ��#7��  �&���Z�
���K)=�Zk�L����S�2�n�3��+Kwpq�*�#�6�Uy��nr|��f�Vyԏf`�   pqM4����, �<{v��痪���x�c�Z������ĭ�'�5"�W���x��Ft�ڥ3�}��I��^O0���i4���    �E3p� �o��1r��V�:�x�-X+�B|����������?�������X]*���^���3 x��4�[   &-�z�G�m �o�3rOf��Rz͸Z��� /�';p�:���GīKwpq�k�qk{�tܷ���[�3��F��    ��9;�h��  �*�:Qu���-U��~���t��\�[������[���[Yjǫw��΀��'17�3 �"��    W 7Q�#"�. �TF��J���{�7��n��/��4����ݜ�S�;��v��GnmDU��)p�������W�Msvb�   pU�Q4g'�+  .�����*^��X��; ��Os�������V�.&��/�݈�N�t
ܷ���[�3��6��I�T   �R�F���  �t�Չj�zD�qyP��~h�͏S���3p.��>���'Jwpq]_��n�t<�O}�^��M� ��q;   @9��(��Kg  \�T��Z�6rp��j��x��\: "§80q��z��#��&"�J�p1��V���k�3�����Ӈ�� |�fpytZ:   `����8��JD��1  �*�*R{9�x�t��Hig�Y������t
���d=z�M�_D�z�.fu���y�t���z    IDAT<��Q���:0�4yv���#   ���a4g�  ���K��#���HU���?��ו� ��L���ΏE�o(���tZU<rk#�̐�#~��{Q7�����    �%O"���3  �D��Qu��L�����fi���;��-�b��L��w��#�c�;��*�x��Ftھ"�-O��w6*��s��   �S38��M� �+�Z��V��D��k�/�>T�Xl���|���?��Ɲ��[��W�n���R�x ��Q����� �9��(�_:   ��#�:Rg�t ��HU+R�y4(�23RT߸������??]�XLK&"���\D|U�.���jl�/�΀�49~��{�s� ">�ݸ   `������  %����nGD*�2R�T��{{�(E������"�_(���l�-������>u�$�Fu� ����^�    �C38�܌Kg  \��^���F����?�}��)�,&���������&�����]����.��+ڊ���l9:=����� �q;   �L�:�Z�� �"��A4���������������O���)�bq���&�1��gZ�U�#�6�ۙ9�q�z�t a�   0��Q4g�� X,����F�ِ����"�ؚWʇpn�����Gķ�����������u����3�b\7�3 ^svb�   0���4�xX: �J�N7�e#���R���>P�X,���r��xmn���J�p~��ڈ͵����>wԏO�uQ����$���1   ��K�h�݈H�" ���F>�W:c��<h��?x�?���]:X�:ܣwڹ�%��g�C�׌ۙI��Q|fߘ�4�v   �9��hǥ+  �\��ii�t��Ki�j-��x�N�t
�܁����c�Kwp~[k˱��Z:ظn��~�8r.]�،�   �O"���3  �\���cG��u�;�GJg �!� f��;������#�U���Y[�ė?��7 3�7>s���� ͸   `�UQ�]�T9�	 ,��y<(�1�r�0��|����V��o.��m{�͈�+a�>�:�*��a��L��Aϸ��fxj�   0ךh�G�U� �⩺����S-E,E��y��J�`����S՟��GJwp>�*�knoF�壟�s��gOKg ,�fx��^�    .[3��̿� �(E���Z*2�R�}���(��7+G���=�ݑ�Jwp>)E�zw#�K^'�����ͧ�#;PL���   H�D{�* ���s#���楤����o~�[Jw ���xY��>��H��;8�����ƪ�K�=9G���cT7�S V��9;.�   �kGٿ� (U��nG�V�i�j��_�y�}�C��d���G�s�~%"6J�p>77����-����N�?*����x���   `!�ڿ ��jE���L,_L���z���*��'���Kڽ���H�Kwp>�K��uJ2��{�x��W:`a��0��QD��)    �ǃȣ~� �"RՎ��f�/.�Z߿����x�`������}����yDx���.��+ڊ��Q������~� ƵW����Q4����9   @���HU�t @y|M�0�za9ǧ���~��[����"�m�=��%��gR�U�knm�3�r��w�=6n(ĸ   ��k�� Xh����f錩�R�������;��b���N?��������yh3:m�̦߾{��Q�����q4}�v    �H3���t @1��i�Z��UU���������~���;?��"ҟ-���K)��nmDw�+"�M'gq��_:`!�f����l�   ����y�egy���s�]��Y�Ui�R��W��Y�L��a��,a���V�m���{:c��nT	am6H�3��тl�D0ƍ��``P-��\n.w?�3��T��*U��y����`��D��y�x<o��3�  �ޕ�d���ye�ŽS?���! 6��fz��;$�݁�ٶePC�R�`]j͎:�; zS�n�b�       �\�Q��c�   D��Ii9vF>��:���� 6�4v ��=W�M�]�Sp���55�)Qt�v'���%e�/�`�yPVg�      g���.+0�  z�))��;-nF~f�C��_�P}�}_��������MMM��L/�݁s7:P���@�`]ܥ�/��� l8�j�R��.     @��v��@  @�2S�?&���PR��#/{��3 t7�H�&߰�j�~?v��@_Q�N�� ��+Zk�cg @�qx��g0      �MhT�X
  z�%J*�b���l�P(��fg9 `�x� ����2�)i,v�M��j�����N��D���K�� Ѓ\Y}I
l�     �z��AV�  �%�,-�;��)�c��������B� ݉�C@�s+��.�]�sSH�Q!�Q���h���j� �I�^��f�      t1o��  =�
%%}ñ3�)I�>����0v���w��M�N��Lo�݁s��i�̈�˅�)���:A�T��N����N=v      6�ZJ�ɸm  �.K��\�ڱSrŤ��=t�~�v蟹Z�9a�/�æg��cn���8w�Li��;X�\��U��B� �9��"o�bg      `���X�]  ]R�*�3r'1ە����@�a�;У���JwI6��fۖAmꋝ�ۃ�W�Z��2 l4o����      �lBG��o.  �]V,˳��Y�\1K~�rŋ�Q������{���Q���n?��fr���N{�{[�ii�; z���
M6i     ���)0�  z�)��J���3�yq����e+��ƀ;Ѓ�g�^'�Wbw�܌��m�`�`ݪkM]\�� =�;M��     ��5��#   �DI���<�i*���o�3 t�
=frv�.�}FR9v��@_Qۧ�ef�S�u��::tlY�K ��x�V�/I�     ��3�L��b�   De��҂�ӈ��+f��|�����|9v����K���h��K����W*��>=�$a�ݩ�:��,0\	 �CG��()�N     @���<tbg   Dg���<;#w�$y������� �pz��R��^�g��&�|fD���5�S��G��jg�S ���L��(9��      �H�P��  ��4 +Tbg䋩b���u�o�c� �7&&�1yݾkM���8{��v��\Lc� ����՚�� �[<(�-��      �h���\�]  �IeXJ��3r�L��F�0v�|cj�[fo�(��4�g�L�ljXC�R�`ݾ7��ŕF� �-��j��s4      "�ڲBY�0�   z�))�坦���Q��v^uom���b� �'6����-i"�����)8{۶jd��xн�W:Y��� ����R��      ��
���  ���J*��,vI���ҏ��~�h� �Ā;��M���ʹ;v���X�&�+�3�u[�����+�3 ������bg       ���Bs5v  @.XZT�7;#W�첤o�C�; �������]m�G�a��1:X��C�3�u�5;:x�*g! l��\��k�3      ��emY�$KM   ��(ɥ��af?ҷ�꣍���J� �§H`�y㾱B���c���V��>="�6"t�V'���%e��v �Hު�[l�     @>y����/^�  HV(K�s�$I&���/��q���c� ��:�T����uY����R��vt�,������) �S��Ph.��       ��g
͕�   ���KI!vF~���P����s}�S ���&4yݾߐ���8;�b��gF�&L��;�K_V���b �H�����      ���vM��bg   �%J*�b|�Qfz�J��G�; �G; ��5}�M?*�-���[��
i��gFU.�8F������V��3 ��x�(�%y�      �x����/�4  ��Y��;��)���?ٿ�%_���۱S �� `���?�H��n��K̴cfX}%��ѽ�/�4�\�� �ŃBmQ��      8{�)�VcW   ��d���9�[�����]�@|����?`�����3�.�R�E��^��MYX�� ��]YmQ�,v	      pμ�&�Z�3   r#)Ji)vFn�i�B�1i��V��� 6��=7���bw��\41���r�`ݖk-}��r� �1���$�v�      `�B�*���   �	SZ�,��������� ��lS�ݼ��N�]`fl@�#����՚m<��w� ��B�*e��      �3t��x�	   I2��%y��$?,��rً����) �`�;�����}B�p�<��>M���� ֭��t���� ��BsE��-      l�Z�g��   �aiQIy(vFn�TR�����<�@�]n���K������/��	~E�jw��YR'�S ��x�.o���       ΫP���b  e�~Y�;#7�l{Z��@i�  �79���&��$�݂��_.j�̈���U�NYp�?RU���N��❖B�;      � N�[��   ?,-�;-�Y>(I2�������_b� �XLZ]j��dZY�k�fb�੕��vmU!��t�\�V��h�N���Y[��(�/�      �y%�㲴;   7<t��{��[6o<�����v� �iK���%����WL]���vt/w��+��F�P__Z     `���   �$YRPR���'�A�O�������0q	t���z������SKӎ�#*xԢ{=trEյf� �-��j��g�K      ��3��j�
  �\�BYV���f���l�=�; l�4v �s3��?%�G��\3�v̌j��;X���_n�� ����KRh�      6N֖J��  �GX�$��,�z�%���w��_������- .<d�.23��IS��
�[��.��`��vt�պNT�3 ��Ɗ�qs      zO�W%��   9bJ�F$c��O\韌���c� ��x�]�-�%]�OmۖA��cg 붰���y���Zk�v-v      �g
-�O   �&I��Ǯ�3mI��I]y=�G�M����.19;�V3�z�<���~M���� ֭���wO��� ���톼�;      �+k�
%Y�(  �#,)H�Ў��vq��������b� �p�Tt��7|��}L�����`YO�� �m��ҡc���	 ̳�B})v      �����*�,v
  @nX�$�N�C�$/�u��j�����- .�$v ��6��}c�ɧ$q�J�V��t��н�m:�p; l4����y       ���Qh�Ů   �SR#���$(���+�~I� O; ���m��\��.�����1="c��T�����U��`cy85�Ζ      �4�Z�g��   �bIAI���0ӄ��S�=W����Kc xrS{��W�~#v�\��j�̨
)�Нꭎ]Vn�����KR�%      �D<�()U$�e
  ��N-��=�$�L��%�bc��w�np~1�����M�w����in�D�ό�\�o�S������:��`��Ɗ�i��       �˃d�,-�.  �+��7E?̒�ŕ�/�r}�}��np��rȡ�׽w4�R���Tb�3��+1܎����?��6�� ��BkMޮ��       rϛ��Љ�  �3��2"�?�/���щ��e[� �O8 w�J��G$�]�'f&m�V�;X��#����`�y�)o���       ��+4�cG   �%%}C�3�dƓ�'�9fb�M���@�L_7�f���O��!��cg ���N���Y� �9���K�<v
      �=<�Y"KY>  �X���9����ʎ������) �9܁�x����R�l����M�Tbg �ׁ�U5Z����P[���      ��򬭤�'9  �
%y�!�l�bI���W}�����[ <3|�rb�u�M<|JR)v�ؖኦF�cg ����Ѫ�MN���se�%�9`      �OP֨Ǝ   �K��ĮȓTI��&w��L� ��@N�J�?����xb�e]<1;X������F;v
 ��P�JY+v      �ݲ��]�]  �;V(Ɋ,�|���f��Ǥ9�c�.�0�����I��݁'6X)�ҩ������:x��v �%4W�F�      `S��C�  ��I����;#7,I^6~Mg.v��Kc �n��=ۂn�T�݂��+t��Q%��N��#��u�� �4����      �&�R�dž�!   9c�B�o��^�w��������np���D49�wP�n��709T*��|fD)���B�@\�����      ����&  <K
��`�<I-)�����.���1�Dd��,�Y�;�x�4ю�<&�}Bp:��p; ��A��$�c�       �Rh,Kbg   �NR��r��0ӄ�'u����- ���@$S�7��\o�݁�K̴cfX}�4v
p�ܥ�/k�ފ� =ʕ�%�b�       ����J�
  �\J+#�1�3�h|b�{bw 87LoLϾ��dv�$N�匙�cfD�}��)�9s��j��p; ���R֌�      l~�#K����   _�dI*�4b��Y����/�F��}ߌ���pL�`��{�$�H��n��]<1��
���>�@|��*��cg       =#4�O�$  �i��'+2��(OT(~x�oyV� g�w`���M����;�x۶j|�/vp�n���Ӑ�Vcg       ��3��J�
  �\J�Ò��3r��F�ʟھ{�1�0�l��={���_�݁Ǜ�hr�S��>�@|:
���      @O�vM��  �q̔�Į�3{�r���� ��s�2}�M?��_I*�n��F˺dr(vp�ܥ�/3� 1yP�-H
�K      ���Y[I�"�b�   �%��A
��)�a��D������k�[ <96�`���h ��"�?vN7T)������9{ds{u�; z�+�/I��      z[�(4�bW   �RR��]ȧI����mύ���1�l o�3�bw�t�墶O�X�.��v ȇ�X���      �o��36�  <����H�|1H���W�e(v
�'ƀ;p�M^��W%�J���TL�}zXI�t;�K��G�� �y�&o�bg       �>Wh,ǎ   �%KK�b�\1�g���ͱ; <1� .����Gd�I*�n���i�]��T*p��%��cU���> 1y��Ш��       p&2Kd)�g  �diI�nH��)�af?ַ�%��~9v��1�\ ���ѾV�}V�%�[�41��:���?t�,��j��p; �䡣P__�       ��Y[I�O2�]  ��L���z�\��~�o�U��8p�wc� x���^�����x��t����˅�)�9yd���d� �rW�W%�K       <����;   �,-Ɋ��3�Ŭli�S��w&v
�G1�\ �����~5vNw�԰�*���9iw��?��p; �@hT���      Ƚ�)o7bW   �RR��>��]��ʟ��l��)�0����?x��?#���ڶeP[��bg ��	:p��F�; z^h��۵�       Βg-%�ʩk�  �(3YZ���Kr���_/���{w� ����7}�����tY�<jz�_ӣ\������?��f;�� =�;-y�;      �9qɃ��,  �3Y�J���LI���]W������f���%��ͤVk�O�scw�QcC}�����G��[�@t:
���       ���uy�;   ���d�H>�'.�ȖW���.z��y2��=����x�pI�L�� �I�����-2� y�P���\       �+�FUr�܂��    IDAT�  �?fJ�FbW䎙�x���mW^���e������]&���x�@_Q�M�,v	p�ꭎYR;c� � 4�\�      t;�Zk�+   r�
%Y�;#w��9�-S7�� z�K �Юk�Wn��K������.�:�4��G�������0� ����v-v      ��!k�
eY  ���P��뒸��4�=�|�����|9v
Ћ�������{%���8��&�|�
������:p��p; �w���j�       �+4���  ��DIy(vE.��������@/bx&g��{�~-vNIӎ�#*x��{,�Z:x��,��* 䁇�B�;      ���
-nm  x"V�Hi9vF���--|jr����NzS��:M]w�N3���8%1ӎ�UJ��)�Y[\m�б��3� ����p;7j       ��7פ���   ȥ�oX��>��]��ʟ��l��%���q��ŁFv��]�S �I�Mk��;8k'�u=tr%v �1B�*e��       .��LI�;   ,�L�3}�؎��x���޻c� ���6�:L/e�U�cw������t��K5�_�� x��\�w�3       \hYSޮǮ   ȥ�4 %�����2~��_;���hj���s�?���)�c��a�����UYX�� x�4�-      �"4W$�3   r)�֩U�8�'��O&~� v	�p���ٛ/��������`Y3c�3���.}�ĊNT� �2�F5v      ����Ԑ;   �Ң��;#��l����Uo��lv�g�����|R�x�H���.����w����ZXi�N �ƕ՗��      � o��V�  �\JJ����3�)��
.����Y�Z
��E�; U����+�@��G�ZZk�N �!4��Ў�       �Ш��T  �ә)�cI��I��붼�mo��lf�����W��}��Ut�b��3�*���A�u���ǖ��`x �&��䭵�       �rI&+�b�   �%)tN���%�Kv^����{�;،�����^���L�GWH�Q�������?R��� �;������       r�[k��9   O�ʃbl�I�!)||�+~�c� �S��S�=W(�KI[b����L;f��W��	�_���;��hq� rǃB}I�63      �+4�cG   �%Yi vFn�4����&w��`�`�a�x
S�S�tU�^g&]:5��r1v
�jͶ�YR�b�  Ǖ՗$�b�       ȓЖ�j�+   r))HI!vF~��p�7�gb�=p^�<��=|�)|F��Dw�Ġ&�+�3���Ro�c��[� �BcY��%  F��
mI5I2�%%g��������5%�oX& �X������_�36��~�J��~;���6� ��)Q:8!{  �䝖B}!vF���y���|w�`�`px�?�����W%M�n�u3c�돝<��զ�{bY�l; 䒷�
�j�  �œ�[X6%K.���$�%�]Z���J�!IZ�aɃ�]V��jAi�^Ȫ#}�k���� ���?�T��N:�QV�'#&��+n�h�y93�4fҘLcrui�d#.3ٰ�c�o �+�)����   ȥP_�w�3�����y��+v
�0��i�\ajr�d�:vJ���%�,�A����ux~5v �Ix�V�-H� `ssi�d�.7�1�N(�{fvL�*�L��|���+�͝�� ��q���ƉN1Y{�y6i�)w�V���t��ɦ]���㱋 �-���
}�3   �ǃ�Փ�B��r�ɠ��nס�-@�c�8��}7�����n�����#2�Rȹ#k:�T�� x2���K��. `��VevD҃���a)��+U��!I/t��ֹV�T  ���+���&��R�m!hZ
�}���%]*�m�"� ��R��E%  ��֚��;#�<����<~��|��"���ӳ7����))������E��:�$���r�:����^�<�< @wH�2=(��ؑ�:li��=ܯ4yh�o~��� �l&w��`(�\li�d�\�,��]��̴M�+ ��e�~%}ñ3   rȕ�-H�;$��çn�l���1=
<l��oޚ��I�����J�T����XHb� O*�Ǘ�\c9" ��  ���q�C&�����w��3�yr�u���  ���\i�Y����g��]��v��s],�B�D ����o����   �㝖B}!vF�y��;w��Ǳ;�nŀ; Iss�ԿM�!�e�SzY1M�sۨ�E�� �:Y���˪59�
 y�YK��(�c�  zG��a�0�C�:`��{'�N�������� �yr��ŉ��;���.�.�|�d����T�� 8��ҁq1V  �xܤ}\W�gn��S�n�'1@��}�g�;cw���L;������W����Ѫ��,v
 �xP�6/9�k �qj����f�M3�F�?b  ��?�n�~N�G-�+�Y�@w���@�  ��	����b��Ss�ɠ��nס�-@�a�=o溽�n_��du$fҎ�UJ�S�'Ukvt�hU�,�N <%WV[��V� @�{�A��b�����j��  @���+M����9���g��/� �L����p5  ��BsU�Z����_�TW�z�K�eIppGO��y�h�W%����.���P_��I��[z�ز���S Ȼ�\���bg  �N��oX���ۿ��_m�������f�2  ����}���ҳ��?��Bx�����c� �����Ů   ��S[ܹY�����w����t��Ӧ���	�����m��h��I-�4���9�� �{�i*�cg  ��˾���%%�ݼ����?�&�� ��{�ܥ�`/�ܟ��?.�g�tI�. �UIߨ���.  �3y��Ш���
��y�w���;�n��;z��u�����$vG/��%�C�3�'ul����l�nࡣ�� )�N �K�����kf��e�/����Gbw  ����s���n��ܟ���0� ���%�K   r'�-HY+vF��7-�\s��;���'M���WX�E�`�^5�_���O!䐻���-�4b�  Ί+[[�B;v  &�U��%ٗ����N�>�� �f7��Ǌ޼*H?���+M�� ��+J�Fbg   �gm��|���~"k��-���N��R��]׾��<T�$=7vK��/�s눒�G�'�Ǘ�\�d) t�Ш���� ���ɒ2}݃��*��_��Wy  ��7���K�n~����ҳM^�� �AR�x�  ��w�� �W���K}~�͛�S`�=g����w����W�����6�B��}ȟv'�౪��N� �Y�v]�Q�� ��\���If_��|�oh�������  �,l{�\+�<d/���K���cw@WJ
J��Q  �3xP�zR{hΆ{�������;�<�Sz���W'������(��v]4�R��v�O�����%�;�� ��CGam^��N �o�<(ӗ/�kI��?�֯�N  �L�^3wi���d/q�J��� Ί���cg   �Nh�ɛ+�3�F��K�}��cw y�U�[fo�(5���-�[zQb���F�_.�Ng��֡c��d�@�pWV���n �&�ɒ��I��J��<��sGcG  ���kn�j��KB�%��?�L��] �O�d`�,�'  ����w�b�t�f�+����)@1���0{K:m'�v饱Sz��t�԰FʱS��YZk��W�� �MB�*��cg  �íᲯ*���랅��-��  ���^���������̮�gϕ�/��iIi�x�
  ���v]�Q���5��{I�|�ɻ�s8v�7��'L��?K>��W]41���J��qNT�:<�; p��R �N&%�&��f��o`��n�mN)  t�+�/�O^����J�Z�/`�;�^��Ȋ�  8S�6/�v쌮�!|i�o��7nm�n�wlz�o�w����4vK/�������iܥ�ͯj~�� �6:
k�y r�%}K�|�e��V�s��{+'�   6��W�8V���]����S�_!�;�9���	ɒ�!   �❖B}!vFw	�����bg y�M��F_���R��5�.��ҋFʺlz8vp�,��j��IQ �:��j�R��. ����%_0�}��/���?�	   g��z��r��=�ԤKb7�F�B���h�  ��	�%y�;��d
����w�?v��cS�ڳ��%����h����gF�$<f��v��G�j���) �u����� �%_P��QP��c�{b7   ?&^��j\+�W��jIC�� �BI*c�B9v  @�����d���jd!�f�����ش�����r��������6�B�u|ȏZ��CG���B� �:x��Ш�� ��f�w��Lw�Н�u�;	   ]`��t|�[�W~�\���w� 6K�LHƣ  �BcYޮ���.�'2���t���Nb�6����GB����J�^SH��6�r1��|_u����(��N �é���x��FrْI���n/�o�{0v   ����fB�W������4�	 �)+()sY  �i<([=)�e����W�'����W>�� �4ܱ�l�G�jk���ٱ[zMb�˷�h��;��պϯ��  ����ڼ:�K �X���>o�;O;|���v�*   lb�lw��J��J�OH��� �RҿE��  �BsU�bn�\��O/���=bz��t���w�\����E�Mkt�;�$�Kߛ_��r=v
 ����ó .�U�>oJ�6��o��9w<v   z��57l���:��Ƥ�R�^ �#)*c   ��l��Y쒮�����]�;�X�d�Mej�M���ӱ;zѶ-���{f�C\[�J�; �x��Ш�� �M�e�͒��mk~ۡ��5b7   g�x��+�ե���n�Y�gb7�ӱ��@�  �\��e:���;��w�C�pǦ1�����}M�x�^3>ԧK&�bg ��V'�б���N� �3ࡣ�6/n\��Ē��u���f����$�  ��2y��x��u&��W��� r)Q:�EJ��!   9�����,Ϲri�ڍ��=ߌ�l4����{�055�yIW�N�5��%m���4A�5�:tlY�,�N <��j|� ψ��f�l��}'M>Y���N   Η�k�pgG�k��j�_j�b�& �����,v  @�x���X��ѕ<��<;����}�5��)��bS���w���cw���RA���*Mx� �����{|E�YD	 �.ԫ�N=v t�5)�Kf����ٹ��A   ��6���J��s���f����	 ��QY�/v  @����ގ�ѕ<��-ܑ�V�c�'zS��z��^����=o��&�uјJ�$v
��K5YX�� 8�]Whp� �^�,�=f�gTX�������E   @,�^3���� ߣ�_)���M z�%J&$�]*  �#��T�/���^�λ��z�[cg �wt�m�p�D'˾.i[�^��i�����q�K�X��j3v
 �<��QX���m �<�*�]�양0����7��   8�ų\i�V~6��(�R����X�_I�  ���jR֊�ѥ,X��K'�z�_�.6��bn��7���~6vI��tjXc����q�,�бe�5�� 6we�y)tb� @.�4o��7%�>y��g���0   p�~d��������N纠ε&��n��ʸ�P��  ���j�3��k5�~�������)��ƀ;���u{]n{cw�����폝�Wout�hU�N�� 8OB�*��cg @�$'$}&M��:���t�,v   �����81��Zwͺ�W�4;	�&��l�   �
�%y�;�k���V��`���r<vp!�)
]i�u{(s���@cC}�tr(vz�J���-+; p�x��Ш�� ��XQ�ܑ�n9���[縧   �PfoI��|s����N惱� l>VTR��  �����3��{�o�����_lf���\sqr)��Iϋ��K��ڹuT�S���udaU�l; l�������@s5]vo�$�������Vc'   ����?�4k+?�{�z�<Tb7�,L��YR�  ���}���w��k�3��QUt��=7�[����%�b�+����&�SУܥ�ͯj~�_l`SqWV��B'v	 Đ��K�%�Z�O.~�\e   ��ȫo+zkO�ߛ�[�L�xfҒ����   ��"��#s������}�;��wt��7�ڂ�QR��W��i�QUJ|w�8:Y�Ǘ�Z�F �l8���X��/���,K���o?�   �S����MwJ�_0�/J~�x�
`���Y��!   ��v-vFwsoZֹ��]7~!v
p�������;Z*��.���-��L�13��J)v
zT�����U�;!v
 �<�v]���b =��[�}"K
[��� v   ���|퍻B��&){����{ t�D���dܚ   I
����b��3v4��/X�ܻ��O��kL��/$����䢉AM�E q,�Zz�����/� �ٜ�nnA� l^�Z�ܦ`�m���|w�    �����A鯺�M>�@w�B���h�  ��`��y����_r�+�/&6������%I���K&F*�h�`���c�5]\�� � \�ڂڱC �sYK�{�`��蓺u��	   ����������kC���ט��	@�%�1Y�;   ��~޸�O/���=�/&6	ܑ{�?�������pi,vK����cfD�,�C�Z\i�N \ ���9%�*��L���۷�]    ����M;�%����?�@NY�t`B��  8�w��O�:o[��7�� �>1!����oL�m�ݱSzE���m�*�I���v'�бe՚l����;M��b� 8_�I�-^�n^���;   @�L�v�ٝ�~I���E�{ ������   ����O�e�ם������)ܑk�{��ͥbw�41��6�J�;=����б�ڝ; p��LYm^r�� ��[Cf��>|�~���x�   xj���[��|����5f*�N�I�Y�#  @b�����/:y�{��x&pGnM��21}I⋾��cfD�����1��M=tbE�9�	 �YV[��V� X'��u:������w�v�������>gf�,�d&3	��e�E�Z��E�UB�~��o��V��ʖ���u�%��m?�E��@2@��E��~j]Z�X�Q ��9���}]�bo�@�Lf�u���/x�29ɼ��u��+
�5    Z�ș���%���A1k����*�c   b���!�WL�<o�맭[���I	M�Wv��g�#���[:�!C}��@��3Y���y� �2�9�ڜu ,Ԭ��>F��x����   �^֞��E
�Q:G
9� 6\��|W�u  @S`��Ҋ!�(ޖ�#q#1Z�hJ��n����k��)��u�U�� !D�d|V��U� �2�iM�T�� ��?���|��ى�>2k]   ���yɇW']�W�^�ú�Js�}�r>c  `�-�K/M?\��CXg ���;�����/�YRb��	r�sȠ����j=Ճ{fT�5�S  �-��)��% ���w�s�S7�k]   �3����S�Կ9J���{ ���[I��
  ������B��_S���/Y� �D+�ʡgo�m���I:κ�d�cTw��X��3�F��7 �	ByJ�Q�� �'Ⴂ����3}�˺!_�.    I:|�'rչ�פQov.<O|��=߳Z.���   ����5B����?�S���e�ʺMۮ��;�;:�sү�T.k��Q��葉YE~����e�ʴu <?�\����щ��m]    �3�!���8*��)Z� X&�+�[+9o]  `.T��e댶�oM�i�    IDAT��g���ɢup�pG��x�o8�&���p��~�]� ,��ݓ��;��A �)bh(�ĩz ��� J�����Go���)   ��r��O��噍J�;��k�= �����s��3   ����y�:���n/ޚ� �up pGSX�����j�H:ں�������� �4衽3�+׭S  +&*�/J��4�y9�JuU����c    `)�q��oSԫ��6#�����L�u  ��P�RlT�3�O�+
�_z�up pGS�t��R|�uG'����C���c�Uj��3�Z=�N ��P�Q����(w��P��ٛ��    ЖV�uŚ$T�षI�X� K�%J��%ǥ�  ��Ŵ�P*Xg�!b�����ɺx*�������~W.�&�>.�L�u�akԕ���l�����(�: ��b��P��� СbT�9w�sn���-;$�/�    :��[_,ޥ�3�bƺ��l�|�*�   siiRJ���'j���o���߭S��a�����]]=?����-��WY��\�u�\a��G&f'��R����u	�N�^9��WO�v�.�    �4x�����.)��)Y� X�;,�d�3   L��}���'���i���0�S��n�+E�κ�2ԧ��^����G
s*̔�S  �RQJk� :���s��yݐ�     �G�0�3ۯM1�yN�4� �3J���H  �t|�|b�o�l��l�CS�if֝{����o����z������3��i�C{g4W�[�  ��bm�:@�Qu'���?1~k��=    �
��������+��2I�u������3   L�FM�\��h_�]^�m�E��a�&�lܾ:��J:̺��e3^��F��[��MU��=�j=�N �iM�� �+J'��i�'�n�?h�    �h���#\��+Ʒ8�A� O����%Y�   S�|A
,�\.�PM�˿d]�2�abݦm��қ�;ڝwNG:���u
��l�����(�: `!�}/"�� ,������$�ţ7�K�9    �=;�[N�z�yR<κ�~$]Jz��+   L�FE�<e�Ѿ��o�������:�E�cŭ�x��D�����F44�c��6U��葉YEf��c��b�b���������;�X�    @;>c��»��ARb���|�*��^�   S�����쾆�={zǇ'�C��ƀ1V���k��s?�t�uK����F�3Іb���Uq��F �d�VR��Xg h'��ɹ����۳���s    �����'(T�/�s���$��x%}Ò�
  �\|?��b�;��]z��Xw���V���g}\r/��hw�]%�8Â�B�C{g45_�N ���p ���K���tm����/���U6C    �
+�s�D��;o8�	!�]�'ȩϺ�$EŐ�gs�!   f��(�˒��^.ι�z���^��k�l�Hlp�
�x����7$y�v�x��RW�?f,�z#�=�*W�� :[T:_�B�:@���sɧ'���uC�f    ���^���uo���V�Z� �|Ϡ\�  @�
�9�ڜuF�K�ӆ��K��:`�+�Wv�d�+�D�vw��*����@���Sݿ{Z�zj� 0*3���u���������_�C    hvѭ=s�Y!�?s.�ĺ�h�+�[+9� ��ҹq��}ٍ�����;�?�Agc�+bݦm����;�ݚ�12`��6S�����5�`� 05�r�:@�Qu��t^WLܜ��u    `�ϼ��r�=
�����LN>��:  ��VF���b�����7�[йpǲ=��SÿI�Z����l��[����ҙ���'{g"'��Št� En� � ��9��m���[�Z�     ��9W��wJz�VY� ����2=�   &bh(�OXgt�(������;й��������ѩ�[�N�Nig�I�:��n�`�g+zxbV̶ $)��� �c���::]Y��X�     ������]�;?��V�8d�t�(�[��Kb  ��w�+Ņ(wnq,�e�t&�x���m�vq�.��hw���iݚ^���=�%힜��  4�X+)T�O�Ԣ�S�ks}�z�����=    ��w��=39������:�����p�  �L1�+�
��!j�)���[/��u
:�X6ï�~|��ߓ��h˨�'���>�D����*�r� �Ͼ+ފ��u
������D����R�    ��������M1���1�9@��!�L�u  ���T�ҚuF��Q&-={��c[*V#�X���k��^`����t��C��x�����;���� �[T:_�B�:@�r���d|��/K.Z�     �@>�G�ͽ*�x�N��ږK�����  @'���By�:�sD��­���:��',��s�}�b�κ��>2�����!��=Ӛ+3� ��P�U�q����W�2����;�c     �k���/�
p.�ĺhG.�+߳�:  �@T:7!E.^)Az��إ�Zw�s0��%7���޹���ƺ����:��A���4DݿkZ�*�� ���iM�T�� �T\���+l��{�5    ��1���s��{�+$%�=@;�CrI�u  ���y��uF爮��~�p[�[�)��cɍ���o]Թ���9�Æ����?�z#���Ӫ��) �f�����H��\��}1Q�c��g�    h]���OIS] ;��|FI��/�  :IJ��%E뒎���ܯN��i��?�p��F6^s�sn̺��2ԧ��^���Z#��]S��^ <V(O+6�� �E��s�Ki�%S����    ���s�8&6*�Q�w���������   Xq�2�X/Ygt�({ql���d��X2������K�S�ӭ[�YOWF����8(�z��wO��p; ���zY��ak������2F}�8�غ    оF^~ٱ!M��69��u��|�\��  t�
��'D���[w��1"�%3z(��������͋	,^����]S���: �lB�t� ��#������/�F�����Ժ    �9V�}�ӳi���Z��c��$�Q�7,�@  @�IK�RZ���,�5�w/ߙ��u
�O6X�6^urt�w$6+,���9:�o��V�6���i5n <N�ك�:��s%���!��ll    XZ��}���݁�s]���|�  :KlTʓ�'J?	��ԩ�S�-hO�����~���oH���)�,��:��!y���3_����JC�N 4�P�S��Yg XY��\V]���p�:    ��6rf~}��PNoV9��u8��!���t  ����RhXgt sa,�u���8h#�}�s�*�vwԺUZ��m��5_���]�
��v ��Ŵ�P*Zg X!1j�ym�udz���     4��mt�P���{�{���J���8  �$�VR��Xgt��;
c����@��e�+��3�]��[�Y.������v �~Št� �Ժ���|����3��9�    h�^����^��H���������   X91*���K:Q�ug^0q���X���0���2�q�W��J�v�t�ak���X��1� x*�<��([g XV�,�3��.��9?a]    �b���_�.T�o��=�=@�r�}�r�� @���z�:�C�{2i��{n�u	��X�u��9;��d���W�t�ZN�c�n <�X�(T��3 ,�˒>�d����=�9     ,��3�G%N��8��uД|VIߐ  �"�u�R�:���/�򯵮@��I�r��O�j�燒�n�����Ç��x���R���w1� ؏�*�/�+ڀ��������̅��/��u     �e�YW�J#V�*��HJ�{�f���Y�  :GZ*Ji�:�c���y��-���@{`��2�iۇ�t�uG�;t�_#�s�h1� �@��!��6U�⩝?d�    �J9�cB���Aw��9��!���  @g�sk����]���.A�c�6��uI���n�v֕Mt��Cr|J� �jC��b� �_�6�X��� �T�k(q7�$w��M���u     V֜y��>����
1���J���x  �Q�ܸ��܊������s��;��-hm�: ��%�5b�}�:��p;�Tm��ln �_L��9� K#��_v]��,��od�    ��&wn�Aal�F��s�s�J�K ����   +��e{�#:ZT8e�M}ʺ���Y,�Ȧk79ſ��hw}=Ys�uZ�� &*�/J�n� E�o�Lr~����f�    @��p�
�^`�X��rI�:  `��T���uE��>I^3~�fM�h�〭=����#I�Y����T��80�z���R=�j ���ʌb�d�࠸�F��c�ۭK     hk�̿<F].���[ 3.QҷV\#  :AZ��ҪuFg�~:�t���o�����:|Oe�n_v��,��8`�F�}�n <�ب1��4��䕅���b�    ���ؙ��0��T��1��{ 1U��ZW   ���k� V7b��K�u
Z�8 �_u�I�{�uG'X���:-��ݿkJ��� ���Beں�"D����
�'�R�e�?X�     к\,�����G��ϓ�ǺXi�^RLk�   ��e�%�\���>w���-�hM�=��Ȧk��Y���U�]z����hi��oה�Նu
 ���b�b�`�4)��V�uŃw��     �Ď�pewQ�?��%NqȺX1.QҷVr��  ���s��9�H��t�p�拿a�������k_'�ʺ�{ؠz���hr!Dݿ{Z�u
 ��z���@Kq%�}6����S�5     ��5/��j�����-����\�W�g�u  ��
���q�
H��CQC���9c]���د����`��7I�ߺ�ݭ�����^�4����h��v ���ByJR�.�T�������|쒯T��N��    �*��Q-�{�='��.�aE�$'o�,�P�K�r>c]  �|�WL�RL�K�8��������6�c�F7m�ZҟZwt�c[��n^ ���(�d��) ����RZ�� �Qr;|�9��K    ���}�I��?,ų���hg.Q�7,9�s  ����-�C3pI�k'n����h<��I�����]��&6�/���n��+�?���,�< &����� �#�}ù�=����պ     <��[_]��S8ͺX..��ϭ��   XFQ�ܸ�u$E�I)wJq��[���qO":�)1ܾ"Fs�	hr��n ���9� O&�{��7Ƕ�&��     4�­[�Z˟�}�)�?d�,��(+6�  �3'�e6�Y8�5r�/J���xJ/�	�۸��t�uG'��e�n��:Ml|��=�%� @ˈ
�))��! ~Yt{��Nz}��?�w�     ��J��yW��n��\Q��vR�u��bZ���$ǌ  hS>Q�3{�,��=��f�r���M�47�P�8������K$��N��������:Mjj�����Xg  ZH��*��3 <�/+�*]�'����u     X�5/y�j��]��!{�{���2=�A�  �e���RZ����D���u=��/��u��x��s�����"�NНMt�ӆ�3Ф�+uݿkZ!F� @��iM�T�� �s�����
�\��u     X�g�J|�L1�Fܚ�6�{V�es�   �"��
�P5���\��i�p~ٺ͉w<ƺWm���臒�8��62�����x�Z�{�Tn ���OH1�. )�}�gܟMܜg�      mjhC�y�����_�n������  �e�ΎK
�!�E�����f���Ā;ct�5/�WXwt�l�u��r|
�Kꍠ{�T��/T ��ӊ6��F��ű���%     `e��������?w��b��U�7$FI  @;
�i�:ߩ7��|��;>��:��[�y�{��/f�}��2܎�IC�{�n ,HlTn�G��
�'��p;     �e��K�\�w'D��\ѺX�PW��YW   ,��Y'��\L˟[����Z���0^�}^�ό������S:A�N8bX��#���Qz`��f�5� @+�A���9���F篕��8����     �ֽ4?�H�a)�^Rb�,���e��3   �\:7.��:����Ή�ϲ�@sa���u�n{W���uG�X�:�Æ��3�d~2>��يu �Ť�I)�Zg )Fw���:��»�[     @sYsV��.��t.�ĺX0�(����.  XR�:�X�ƚf�3=o����Zw�y0������Y��!�Nq��k���Xg���,i��u ���ZI���h`����һ�c�ۭK     @s[{f��1ƏK�8�`!\�G>7h�  ��B�t~ܺO��ٴ����/x�:́�P=�\!��WL.�p;cz��p; `�bh(Tg�3�N3��+��x��     �@L���Rػ�Q��(W��TlT�e�  ���)鲮��a��k)EwC�;�ȫ�=݅�o��Nq�U���@�(U���)��S  -%*�/J�nt�U���e�˽w����u     hMg��v5�9����)k�<5/�7$�Y�  �G��*��x�g�9�㒫�;`�����k�.�7�K:E&�:�a9>y�To����`� h1�:�X��� :��)Qr�ޱK�.     �a���)i]����[���J���x	  h1*����Vs��Iw�{o|��v8�@:�Ȧk79ſ���$���:d��:M ���vM�Te�. `abZW(�3��眿Oޝ7q˖��[     @{Z�a��Q�����[��q]�����   K&��e�<��V�����s
��%��q��/u�\�+���[:��F�I�u��O�g5[�Yg  ZM�
�I)�,?#��<�?K_����k     @�*����˧��޺/K�y�����'���.9ψ	  h�3���b8�ow�|�����)���5�i����a�N���KO_��:M`�dI�'�3  -(Tf�%��]Ey��ȾsⶋvY�     ��2x��L\�c
�U�{|4#�(���  @;�J�&��Z���8_Vw�Y�x?K�:�h��+G���#�i����������nj�����Xg  ZPlT�mo�����˼c|��_�n     �m茭/s.~Z
ϰn~������3   ��Z��|��{�su�&N"t ��v��2�����I�r�w�R����  ��*��Z���K.�x�Ng�     4��[n+�}��(^����~QlTk� ���9�<��x�P�ދ�3`���s�9!����2�-�d���΀�FtϣS��9L X�P�RlT�3�v�:�>_w=��qW#     ���~��#W�<��&I�u�����K��!   -���B�:���%���6Ϻ+��3�iۘ�3�;:ͱ��Qo7g
:���5S�Yg  ZP��*��@ۈ������7�k�     p �6�礫��,�@��%}Ò��%   %T�ks�x*>���a�N��o�[�`���AF7]�21ܾ⺳	��nWq��v ��T�2k]��(��K��o��:��     �������\=G.��(W��S�ʌu  �As����8i����Yg`e���S�0��w9�d��i���`�u�L�W��^�  '-��CR�A��!�s�҅7}�#     ����p�H=�>.��YhS�{@���:  ࠤ�)���E�p=ϛ��=߱N��`��C�n��O��6�Nt�ӆԝM�3`�RKuJC�N ��P�W�2���_]&����     ���q��%w�s:պ�����%Y�  �E���2w_w��+': S�`�9�p��W$�o��i�z�lo�g��    IDAT�P!Dݿ{Z�F�N ����+��@ˊrS���8��-��_�˺     `�������׾���G��(���z��Йb�&��I���  �59�(�K�8 a$7�H�w�k�%X~\Y�|O�bɭ���Dkx�ԩ~:>�J�a� hIQ�2#�@��sA�9��g��$     о��0�s�vɝ,�,^*�BL��Y�  Z�O$ύ4-#T/\�{�8�:ˏ#�mn�ƫ�]r�8��✓N:r��ǬӌO��ha�: ТBe����"��]�ɱ�ߴn     �0r�egD�W���nA�q��]}�   �j��Y�(��V������,6����2��&�{�n�@�vn ,Nl�n���%N�U��    @'�yɭ}:Q.�Pr�hĊ��Y�F�:  `Q|�˖��Y��wYg`y1}��F6^s�s�;� ���G4<�|�$Q?~��z��a �E�A�|A��u	�B�-J�\���G�K      ����<2q��)��a݂�%}ÒcD  ��t� ��uXR�I���[�w�u	�Om��L��ͬ�uY'`��t|��v �����������(����ֳn     x���?Tؑ��}�):�����*-O[W   ,�˲̶���kۭ+�|~nS#�9C.�غ�S��d�����$��eM�W�3  -*�ˊ��u���kH����;�8���:     �ٍ��rCR������{�,���P���   X0��N�B�ڋ���o����p�X������t�uJ�:t�_#�s�X!�j]�>:��K  -)���:�� ���k��������K      Z����ω>nw��Y����ܐ\�[� @kI�R�[g`��SI��	�7��n�,-VL����F_�p��U�<�w�4D=�w��v ����i1��G���%�*�m~>��      �W�-���sݳ��y��{��BeJ
�u  ���Ž��cij�u����Qo�|O�T���#�[:U�;��[c�����M�W�3  -*�����@s�x��2�3�i{     �%����.�6�Y�-hc>��wXr��  ��CCa~�:��z^=����u	�Omft����#��l��>�[�k��0>]֣�9� @���`\��5 �/��O���O�m�ٺ     �����uc⧝�!�-hO.�#���   8`����X(����������u
�������O����n���:+�TmhW��v �bE��n~It�̕����3�     ���wl��gKϐ�ՒR���ب(T�^  ���N�b�t��\��:K��mdtӶ�Jz�uG'�&^'9l��eB�=�N�R� `qBuV�6o�4�m��G�c�}Ϻ     �m�?��p��N�nA��A��  @K�i]�T�����$��ޛ�w�u�m�Ѝۏh��ǒx"4�f�GG�Xg`�=R���t�: ТbZS(q#�s~&����s땒�Z      K�]Cs����>��w�XB^�oH�g�C   �R:?!���"����'�;�Ϊu����h��b���@��:�l�\c� �x1*���+����#�:����O3�     �n�׊c�-N�Ӣ�7�s�N�ByJ��:  �)q�L늡~�df��<6�����l;E��',�;��ae~�*Q?~��z��. ��	�i�:��(7᝿xb���-      x2ѭ=��?
!�s�ںm"�RһF��  �fӺB�`��E��ה�������к��$npi�B�,��vgnos��2� X�ب2�HrQ7t��D��     ���;�l������A�Hk
��
  ��rIVr�u����Ci�uGb[���k~�9����֭���5}�X&�ي~:>k� hU1(����Ut�������-[��:      7�!����	'[������.�_  �+Tf�%���������Zw`qX7��s�n�>�.�,�Z#��u �������dQ�!4r�1�     к
c���g��r��-h}�:�بZg   <)��N�AJk�O��x�u��-ld�ug:����tґk��D���vMi�\��  ��X/+T��3 Q���Ͼun�n     ��ސ���x�S<Ժ�������u  ��Jg�%�̮�ez��p�o���±��eE�b`{{���u1�ަƧ�� /�
�Y�
�B*��z�W��p;     @�)��oL����JrL�`��Bi�P @�rr�.��F�uk_�߶���1�ۢ֝{�c�c݁}����u�X���b�N ����4)�5�`�����a���b]     ��7�!�;�q�\<ƺ-*�RһF��  �fÍ�m�e\8|�d]�V6ݶ6����31ƭ�����LkG��2� X�P+1܎��j���>z*��      ��0��߹�էH�jI�uZPZS(38  ���t['`)��3����u��-hݦk�宷��>�9=�r|��Ja����g�3  -*�u�RQ��1~���X�-�-�      �93�[!�ϲ��Ჽ�=��3   #�/H���-�'e��2~���Z������������K�;�s�=���L���0g� hYQ�2#����kH��B�?��v      ����g�ܯ�ܱ@�^R��[g   <[��DHs1V�[g��1��bF7n;_N���ϭ_ӧukz�3���3����u �E�ʌb�d�,����8>v���[      �|�n���cL?�6w,�����Xg   H����XN.���������%xjlpo!#�����;�X}=Y�,��l��v ���F��v���mm/�g3�     �'31��kls�b�ʴb�f�   IrIVr�ڶ�(��O�{�G��K���Ե��I���9���u�H���ȕw �E�A�2m],3�#e�
c�w�<�0     `����ra,�N���(�{�{�*�BeJ14�C   $I.�m��%C���L����Sc��E���k%w�u+ו���:K���i��  ��P��"K�Ц~���Я�
��e�     ��2�3�u��cAbP(MJ��o �=�0��Vj�?~�ǎ�����z�E4��$�ʺ����G�]̕뚚�Zg  ZT��e�`Y���c�M�^�]�      ���o8�,�k7\������c����b��4��wh���   F�mpw��u
��S��Z�JI/�n��c�{X���H�m�x�\w�:K F��Y� @�
���@��r�����~m�6��     �4&�6-7��9��控�J�Sb�  �rNJ�l'�Q������+�;��poI��I9�<^����`�TI�:��  ��V�%qE*ڍ�۹䷊;��;�׭k      �^���rag��N�����A�K�
��
  ���mqG��J�O����X���1���־r�!Q�-�x��;�t%�8H�F�ީ�u �E�ڼ�֬3�%�s�3ewja����     @{����������Xэ����Bu�:  t0��Ph9W�{�u������n��)�ͺ�ן���C�3p��=���� ���i]�T߹�]D%?��wn�'�      t��g�ω!n��z�4/߳Z.���   *��bj����J�o��=7�����ܛء�!�?����ue�p���� )*Tf�p;�D��_��3n     ��������}婢'*3���  6\��:K-�=iy���x<ܛXçI�^�&���Z'� ��H�+�  �*�R�[g K���$���3���X~ƺ      �mz������I�Q���A3�
�)Ŕw�  `幄q�v���k_�[w�poR����#�F�<��n6�����%��: Ђb��X/Yg K�ݒI���[.��u	      ��
c��rI��Q���ByR14�C  @�a�{��R�z�1��Ca��I���,��T❺��u���*[g  ZQ
�i�
� ���
c[��s{~�u      �D
�\�Hq,�R�?�4o݃&�BiR
�u	  �$�K�Ÿ�(���OgJ����1�ބF��~t�{�u�\O�I��]�9��3  -(Tf���r�2���eN����%      ���عe���N����nA�������  �����]��z���Of݁}poF1�,�	�&����U��55W��  ��X/+6*��"�r�?�0��ES;/~Ⱥ      X��.���\� :�5�լ{�DBCiiRb�  X!.À{ۊi�+W>n��}�u k�U��p�poj��kdu�:�p�S��ԭ3  �&�J�����������7_�C�      �`�l��� �EI'X���$]Jrk$�  Xf1(��k]���|�����+��W�N��&�2!/�ۛ^O�[��\��v �"D��i1܎�J��!7���     �.��.�^��Y��Jr���>iMiyJ�� �2s^�Y�
,�\�6�99i�@Y���?��	G�+Ï����_Uo�� �0�:�X��� $:����Tܹ埬[      ��v�ֳc�����-h.��ϭ��   m�9�v��2}0q���ƺ��1��DR.?���x�p{�.3� X���y(E�q�})��L��     ��&ƶ��;5*�ͺ�!6�
��  ��\�e��ec���l��ۺ��%��g�Uۏ�>n[��^�+��U=�X�4D=�wF���  �ByR��B˘�1�Ӊ[�V��b      ���=wΕ��}���nI�#)k�c�.Ir�  ��p�+�J�XN1��eU-����[�t*�P7�$I/?����Ź�V�w��40� X�P��B�:8 Q��i���ߺ��-      ����[�;�N�ܷ�[`/��j��  �]9'%��lw�Q����k�[wt*����ۏ��j���,���.[g  ZLlT������jQ���s�[S����      ,M���]ػ�ף����&.Vgy�  ��K�-���F_�L_n�ѩ�u �u��}.Jo����9r�*�u[g� =R�c� �0!UZ*H1X� ���=J���m�oY�       �f���o�Q���n�-����Xg  �6ӺB�`����4����x�X�t6�[��G��8p]6���Z#�0�p; `!���4��hv1�_��[u*��      �ߙ�z��i�%7X��V(O+�5�  �f\�#� �I�W?e�щ�t�.s���u\w��V�{r^1ZW  ZI��K��F�r�蒍ű�[��|N�      �1uc~jb�Mr����u�D�ҔbZ�  m�II�:+ ���}��ϱ��4�z�5O���;p��xg��P�����Xg  ZHLk��9��IE�o�_��=Jһ�����Tu�=�If&٨���o��!@4�8	!r[n��LWѳ�+��@�U�(A&�=D����芈@��LwU������}���	�LwW��.��99�9��;��Lwէ����ק��ػ      &���/������-�Z�Tx�  �J��	�&���W��1�M���Q9eo���pCd���Ccv���v ������xV�����=c�p�.�      `���bm�ާY��.)z���%�f��;  �Pb�<.�螹����zw�NQ;9������I[�[p�v�آǞv�wE�H��Wk� ',�dO���1�;�M\U?r��x�       �b��מ�,�����n��PR�}�BV�.  �Β�ʬw6K61'v~�a�;ep��I9�7�q�Й,�%3�� X�[��1��-y��D��      @o��L͔&'Д��wXTj�K�C�  `�B&e\q)�SN�k�3����NS̿$i�w��Swj��m�xEL����J,� '�R�ԨKJ�)�7j�~�:3�[�!      ���{���6�;d�7��M(���)+y�  �!��K��靁���c�����ڻ�SF�=��ĸ}(q�}��-�� N�)�Ÿ��,|Z�ē�      ��:=uS&=M>�݂MfQ�Y�;  ؐP��X�bk�i^�1X�n��ܰO
?�݁��`�>�b2ՖZ� �!���Rʽ3��B�tc}WxR�����      ���t�����'*�~߻�̢bk^2��  �ub�>~��U�_�k��1����&���A��݁�)�x4� �-��� �Ί���0J�ߪG�;�      ��c���!�ŧ^xݭ��
i�w6I*��*m�#�� ��	Yy�{>07>,��n�m�.�Ne|g���^�ۻ2�g�;�~%�d��T�z; �DXRj/zW �$��7��      ��v������K��[��R���;  X�P��N�&��{������Q�Zwe[�?m���O��)�
<��fGy�� �G[��@�A-do��Ω�T���      �u��~�6{��,do�/(�F�  `�J��tI�Yy�w�(c��I�<��-K��_�t�w�g�DI���N������Zi�� ���Yg�;c/�'�~�vt��%       ��*�Mf����-�$�I����  ����+5k��tA��ݗ�~�u�]2���I�v�_&��Cm�̗ˠju�� �Ge1�uV�30�����1��v      `8T�+�$O�e�݂M���y�̻  �P*�{��ȔR�m:�R�.E,v7Á�$��;S.��2���-� �����Z�ċ�p-do��~�ح�Y�       'n�h��ڮ�=�B�v)$�lF�  `M���qGVt�ܻ{�˽;F��x�-��;�1{woӷ���;��_�)�� ��ւ�h{g`L��=Y��d���'�[       l̾�?/Y�{��y�`�����d1�  �&�e9�Z�Q(M�7��=�_��n%���;&�w�
l\9��e՗ی� �(u���Ɣݚ��1n      F�����!m�!)��l��Ql�X  ��B6� '���l��;F1�Ӯx�s��w6�Swj��m�x��}��N�3  �bW�9/^x�f3���tp~��ۼ[       ����Nm|�Wd���J�9�Pުl�n1�  �b�Ԭyg�K�X,N>�;?�y�Q�I�>3�7y7�7��T�r�˸ ��,)�Ÿ���.����      ����X����Y�BY���AY��;  xD!+�Í1�w�W����>�w�;�!�l��F�����.��  ,�%�P�lᖴ%���t�/�K       �_���ǂM>���w�,v� ������+�)v�+o��1*��QP������ɣ�[]� ��J�)v�30^�)��6S�h�Õ�       ����_��>Sy�)�N
ɻ}��  <�Pb�>�R��Ӛ��;cT0p��W��$��wz���`�]h�x�  �,ve����p_�Jϩ�T���w(      �X
V��Le�|�)T�k�G��؜oX �o�wt����������Ĕ�,�E��_.�"/�V�� x��Z��'f�����G�>�      �������\~��ɻ}��-F�  ��Bi�;ެت��A�Q�b�N;p�w�e��-.���RK�
  ��[�E����kg��=��_9�      `p,>����gIٍ�xcsT1r  2�_���o<ƻc�1p���K�Y#&c�>b2ՖZ� ��:+R�zg`�4����L�jU*ɻ      � ��o浙��!�^(�%��	#w  ��B�2��cϊ-Y�5�1���طx�)�^�݁�c�>f���  dEG�mxg`,d�`����#��z�       |�#�?4��J�w��I�*6�q  H��;$)�x��7|�w�0c��c]uV���^Lܽ�ERu��� �IQ���]��g!���v���+wy�       ���g��<�	
���[�')Wl�3r  RV�.�@���a�b�����mm6[_�t�wz)�    IDATs�w�ػ����w �72�F]J�wF���J?];r�7�       l���}����
��݂>�&TھG
ܛ `\Y��HV�rԶ=�_����w�0�;�j��/�����v�"��̸ �@��̸}�}&d[���      @/T��n�D��p�w��K�   +{`PXQ
ݕ�3��^�T2�^�<��ݽ��yW  ��-Y����(�?.�gU����       ��v��?X���0�݂>`� �XY�;�b������zw#�=���N{�L�ٻ��w_�v��F�; 0@,�J�%��(S�Z(��6=��n}Cû      ������3��J��J��=�1F�  ���I���,f����:0p�����	,�ݘIwWW�3  �ĒRkA��@?��2�~�>=��       �.Xmf�R��BS�zנ�R�ج3r `���:�݋N;p�xw��z`߁��t)<ջEե����; 00����٠B�wab��3���;      ���=�KK�d
�ϻ=�
F�  ����]�Ab1��!�a���B\oqf\��PĤم�w `�����r��Y�jM�S��/��      `�,��yR+<U!{�wz,����8� ����;��\�����w�0�h��x����ߐ�[�_����0v�:��f��� �U�ېu�=��+j�So՝�qB      ���;o+Z����[���ǂ�GT�nB����(��(nQ 0�,�R�x��e�����O��wɰ���Bx��uyp�|���� ����+�,{g`Ԙ�H��Z���}�       ���t�=�P�QS����ĢR�.c� ���mx�w�8������1,�*ڀ�ܰO�yw`s���}�1�k�� ���T(��30bL٭Eiۓ积�W�       x�ٙC=�����nAYRj�3r `���X.:�k�+��Ha�5��zw`s0o�<���c��  KJ�yI����������y�G�<�       �ح�����=�B�v)�B��8�އ]�  �/��;���O�r����1��ә�߰E���������Xht4����  Sl-H�C0"L�j�.��T���7w       �͗��t�!�^$<{d��^t�C  @?0p����̊�/yw�봸�t��ӽ;�y����n�t�ܲw `@����^�����*�U����       kU�>��Hg���-�Sj-�r� 0z����Y��l�7�'�A�W�:�^�݀�UD���Of�]�K�\� HJ�Y�������4k�ٙ�_�.      ������R�����-�Sj/�  ���x$VlQ��F�AǗ�:�v��ϲ`��������N��;�xg��{��.4�3  ��R{�;�!����g*S�!       �;N9��J�]#�GDزK���  ��JͺwY6ќؾ����|��wʠ��uH�~޻�//���/K�.�v �$Ɋ�v�),�L�g�      `���T��R�
I��5��,+uV�3   �R�=�6^�1���Ѿ���t�w6_���	#�ݍ�kv�; 0 ,�J���������G�;�       �2w���rv�)��wzú+J>�  ���E�=n��1���Q(�׊_����2p�"&}�آb2� �3K�Rk^&`�,�H��Y�3��       �V=\����ؤ?�nAoX����H  Í�N@�w�;�?�1�����|�;N����UI;�[��&J���zg�3�K�-h��{�  �Y*����a2lH4eo��T��C       `�Y8�k�G����d$��6e�N�8 >Vt��Y�&�;�}����/k{�.����ĖW�q���cR^$��
�v ��"�vl���J�0n      0��է+oTVz����k�qV��Z��,  È?�qb,�{��՗xw"�'��JYA?�_+mٽp�|C�%^S��gI�Yg܎���,������a�       �V;2��a�W�[�qV����H  Ã?��)uߠJ�=���r���?�RI���V�;a��-�tl�� �Ƹ=`!;&[O�N���-       0(����D̞h��ڻ=;��y�x�<  C��;����w���΋�;��~޻���oHm��{j+�  o���R*�K0�L!{[}z�yՏ�m�;       ͱ[+���{�)���nA���{+�� 
Ɵ�XSjw~ѻb��a���w��̲Oyw`0�y��ڱu�;c�,4:�kv������q{�]�����e��9�~�       �\p�Jz{��aJʶ�Q���%  ����,ozg`�d�v��]�W�%���' ��j���r�;a�ԗی� ����>��ٌ�      ��է���&�3��w6ȢR�.��� �@�;�,�:�7{W��+o�+�
���FG1��>Qs�-}un�q; �;��ذ�S*M<�~���z�       ������d�IR��l�%�漬�z�  ��a)z'`Y�w�e��>�A���Q�_%i�wGL��b�;c(�o�ڊw ��%�f�q;�/dأSή�r�׼S       `X-��i���Q�lTRj��r�@ �@2�X�!/��;cPv�����z���z�`�����}̩*e|	=3������0 c/E�ּ�
��h��Z��Ly�       ��p���V��A�za�.e�;�3  ���W�yW`HYV�f��|G���o\p�C�b1n�C��tl��1��"��.0n ��ۛu��X+Yi���      �ׂ�g*S*e/U�x|���βR�'� 0(��6 �bR���;�G`���n���[li��{g�F;��_�W�ͯ �����<v��E�)s���w       ���-�߳�=[
�y�`c����^��   G �a���{�o�������a�~�=�ҹ�lw�-)&��ե��x��S  �,�۱�_�){r}��Y�       u����6������{�`c,o*�$�a  ��%�ؠ���R�����?���I
�ly�t�E�1�1�+ǖ���l|  �Y*���۱>!{Om�㞽��J�;       �E�c�r�]���t�w6Ɗ�bs^�y �#.����ϪR�7�p���8yrr�ݒvx�`8��}R�=m�}E-4:�ZuEW� �,�J�y��sk-��T?R���!       0�N���7��/K6�c���M��}��� �f�+sD�w��؇^��/|'��LN�L�۱Kͮ�2�46��W/�/�+ǖ� $1n�X����<��       �6=�����X!ky�`R�بɸ  ��J�q;z�;��yWxb��M,��OyW`�,6:���u���*%��bK�����F�; 0 ,v���۱v&ݕ�윹���       ���-S�R�#��^�l�E��,��%  ���E/Y̟���;��ᅁ������%}�w�S�[����k~e���fR}����]�=��1�T xtV��q;�*�c)dO��>���%       ��>�V�Y2��0���{׻ ��`��;zȒR����^�?H�����Lw�.�{����}�k���ܲ��" ��h+��%��'�Q�>P�Ξ����       xh�+w�������-؈�:r/��!  �<+�Pz�ȯ��K�y�w���w� 9��M�I�n��@^$՗��I�&���U�j�m�5���R[Ed� x ��J�E1n����֧+?����c        ������n���}�_n���{�~��Cyҹ �eI�Y����I��l~���]�نgq�	�,�J���c��m���y�qς�W:��6;��[ֿ�U�=�usvg �o�:n_�v�M�
�tU}��F�       �Z�OWި��3fʽk�~�]Qj/��x  �=���oR��z�M���1��έ�w���$��N�hʋ��FGե�Z�B�L�R�R\���Bե��V]��BK�n��� ����Yg�;��¬�tAmfj�;       �>��?���|��X���ݻ�r)E��)��  %�7�Txg`Yܹ��}��[?흲��N��}W��@0}л�gۖ��o���ɒ�o)k�DYY�F�fR�[����h�Zi�*b���/ ��I�Yw�;C'�lQ.=w���/{�        6n�y����E���n��&U�v�2�  FB\���-�#�&��z�5����L܏���W�g{w ��e���rI�r��R�r)�dy�?C
A�BP���L1��UĤ"&�ER;/�ɣ:ݨd�g �]j/��w�N�eK9\q��
��       �����މ��4Ȟ�݂%e��(de�  ��ŮR�����s��fo����.�,�%��ߝY�9��  � ��Z�-��k3׾V
|�       Fс���O�^蝂��m'+�&�K  Z�f���~�����Iʔ�Z��  �L����k-�__���j��       0�n�tkӕ�Jo�B���:YRj���w	  C�
�E��ؽ�K޽߻c������/}�V�^��  0P,)����.�P	Me�ק��w	       `sԦ�~U^",���)�d].� �VVt%�~�`�DJK����,c?po���K:ջ  ``XRl�K��]��rL)<�v���x�        6W�h��!��3��݂�K�%���w  C��w�H��W�R���X�M>�^�   00RTlԤ�{�`�X�\����*�       �Q�9�Y��4I_�n��Y�Tj-H2�  �%Y�Cl��b񘽟�q�w�f���+���
z�w  � ��+6�E���Tl;k�h�N�       ����[�0��O����n��Y�^}گ%�  Z�[�Ca�\&���zWl���+駼   �]��<�v�M(�~�����M��)       ��p��[�v��L)�c�l@�FJ�w �ñ����|��~�;���o%� /���A�w%m�n  �dyK��(>U�5�Jv�v������8�       x��;o+Zw|��m��W'�S�{�N�dE[�4����� ��dEW�7�30�,KY�m}���.駱���e��N��   ���X����JW�>v��x�        Y������k̔{�`�,)5�eEǻ �������'��ez�M��4�w3�ܻ  �Sj/�:��.s��t?�       ���ԻK��|)[�n�z%�ּRg�; ��`��"��K�}{g�»���r�~���~Igyw   �0�ւ,oz�`����r����k��;       0\�f�f2�sM����uW��K��� �qg��c 䝟�N觱�'��   .,)6�eEۻC%�S�<qα#o��w	       `8��\�ϊgI�3�-X?˛��yɒw
  >Rds��`��}�%�����2v�3ϿaK0�I�  �M��b�.Ůw	�JvxW+�=��_:�]       n�[��j��1���݂�]�f]�
�  6]꬈��` XR�#{�}��˻J�J:ջ  `3Y*V��Ј5!���]|�m>~       艅W��>K�����
�f]�a% ��TȊ�w�u)^q��7l��臲w�f3�^���g  ������Z�ģ"q��B����Ե��N       ��O�f^����'�����%�漲�')Ll� �דּ� <P��Y�,.���^����;��   �źM�ּ��D�B7��ק���n       ��`���7&e?')z�`�L����Y� ��,沂��c ��+��a��)�^�1�{  �+���:K�&�-J�ys�S��N       �����;C�]*��݂��nC�9/�y�  ������R���/~�c�;zm|���V�Az�w  @ߙ)�dyӻC��.M���ʭ�-       ��R=R�hI�7��݂��f]J� ��[Rʽ3��f1˭3rW��f�~ھ�H:û  ��,)6�<k�}>Y8g���O{�        ���̡���֧��[�)_}�*2 �KJ�e�
����U���&|��fI
z�w  @?Y�5>5�51e�謅��;�[        �:��/Lj�YR�G�l�E%2 FD�H��3�G��o���;���Kc1p�������   �bE[�Y��G>�ąP���N=k�Õ�        $龙��e��LS�g�-�Sj-(u�!  ��Ů,ozg '�;�W{W��X�C*�DRٻ  ���Tj-H2���{�Ӈ��͕�w        �h��J}���W���݂���2�c ���R{ɻ8a��sϸ���2�,؋�   zϔڋJ~���t�:}�+����       ��t��6]y�I�{�`c�h+6�%K�)  ���]�R���`�D�U�wG����}���<�,��  ����ب��w	����L�+�3S�        
����Pz�XG��Ul�d1�. �QY�e݆w�fV��{7������ �H��+6jR�@�I#˲K�f*��       �Z�OO�]��2S�z�`,*5벼�] ��3Sj-xW ���=��_�wF/�����/}�VI/��   ��[Jͺd�;C����G�ӕ[�[        X��-��+g�IZ�n�F�R{A��$ɼc  �&���&C,)���]�#=po��K:ٻ  `�L����^/�a-L�n)�H}��w�-        l��_�X(g�J:朂���؜�,y�  �,oɊ�w�!����	遻��Ļ  `�,)6�e�����Vg�g*��.       ���+���&�1˾�݂�]�FM�
�  d�Pj����=uou�|ف���x���xw   l��\�Q�b�;C�,�۸Eg�����       @/��r������쟽[�A�uY��. �33�֢$�,��`yg�����=��%��;   ���Rs^�蝂!c!ݾ�g/|����       @?��2kҹRv�w6*)��:<� �#���{g ����i�w�F���]�^�   �>��YVj/�Oc���ԟ.���׵�K        ��Lei�N9O�>�݂���RkA2�N ���Y�I"=Vl-uxgl�H�O{�;�����   X3K��yY��]��cR魵�k_�J�OF        ��3WwjO�e!��z�`�h+6k�Tx�  ƀmY�'�`D��E�	1�w��%�   ke��بI�띂�-�^_����;       �MW������4e�y��R�ԨsM �Ws�֒w�7�����m��5r��;��I�.��   X��m(5�E�3�e��OO�û        O��ʔ�����N�^Rj-(u�� ��Z���#�RV�+�#7p�ͪϗt�w  �	��؜�u��K0��V�J�V~׻       �AP�>�k�e���»gݕ���w
 `T�)�8@���R����5r�`�  `�X�5)v�S0��%������G�K        $sG�~;d�)4�[�qV��u)1D l�)�楔{� �#���w����X������"�<�  �GcݦR��'��^s!�Ϫ��s�        Qu��o�e����K�b�&+��% ��eJ�E)�g	�IRj�^�]�#5p���&�;   �����:K�x�"���V6�#�#�ʻ       �AV;:��L�\Y��nAXRjՕ:+�% �!�ZK���l�B����V#5p�t�w   �ñx�e��w
�U�nOa��#��;       �a07s�?�,�c�W�[��]Ql�K��S  C"���j`|������i�k52��t�;�]���   %uJͺ�
�)ٿ�=}a�^�       `�ӕ/H��e�s�-��Ql�d1�.	��:    IDAT ��^��M���)��Cw@|d]%i�N� �gI�9/�,K2�)��7���#�n��U        ֡>S��;Α�Oy��G,*5�J݆w	 `@1nV���R���P�>���n   �FV�U)v�S0�,��'�ó�?��E�        ����J5L4�)e�y��WL�YVj-H��c  �q;�u��{�e�9�k1�}/x�K�~�   I��R{�Ұq��~����;o���S        Տ�my�N9�BvĻ�cE[�Y���; 0 R{�q;�`E�B��{H�*�   I�T��x�Jؠ�߮�z�*>%       @�1su���q�
�݂J�R�&�[�%  7��Z��ࡤt�|��q���^�dRx�w  �u�J���r�����t�R0�        F�͗��L兦�7�S�K��^Tj/J��, 0V����q;�P,��N-��#�'j��}v��$}�w  c���J�%I�P�1Yv�6S��;       ���>Sy�I�{���,o)6�R��) ��`i�����.Z(�z7����[Wy7  ��eyK�Q�$�BT�~�v����!        ����u�L�u�豔+6k���� `��x�CM�w	0�,���Jٻ�D����/}�V�]��  Ɛ%�����&�;E��U����)        ���Le*��7����KJ�y�6Ob�Qd1?>n/�S��`�)�O��,�1��f�}����;  �x��j�m��S'+�������w
        �l~���C(�FR�nAoY�Tl�s�
 F�m�f]2���"����'b����  `�p�=��B(������K        �T�>��,�_(Sǻ=�ǏX� ��u�J��t`킊���K��fh�g<���t�w  \mG�eK!Vg�{�        ����>�A�KW�o�KJ�y���E�02���Rg�;Z���}񮳽;����m鹒vzw  ���v�I5%=�zd��-        ���n��S˲�daŻ�gyS�Q���; p�,)6�ey˻z)�^���h�v�̮�n   ����
W��ss���h�c���        �>=�g�ҏ�4�݂>H�R��P ���\�Q�b�;���;�����{�o�ʶv�I���  F��b����`�3髥�mϚ����n        'f���Rv4��z��?By���'Iaho��Ȳ����y� #$�<���}�u��]�p��l[�"1n  �f��YQ�S�����ɲg0n       `�T�\�)��3�p�w�Ê�b�&�=B  ��^Rj/�q;�k��ڗ{W<������  `�X�QlTe�����6�s�V��        k7��lb�9&}ջ}bQ�Y�J0  K�b�.˛�)��
E~�w�#	�ku�U7�T���$m�n  # E�β�h{�`de�͂�=7]�        C��;�������-�lB�m'KYɻ Ǝ���6J�)���,������_{�w�C��n�R1n  fJ��ի���7�g�Q�d�       �h8v��_��tI�{���R�ب�r�G�Mc��^Rj/�q;�R(5��+��܃���  `�Y쮾 �]�D���OOh�Y�n��z�        �ީ�T�Vi�R�y��SRj/(�%�=E �'K�b�.˛�)�XIJ��nx8�;`-v��]{��OҤw  B)*u��؎����S����?��E�        ���W�;��'B��nA�eee[w+�&�K `�nC��@!�"��߲��_Q�Ny����>Y�Kĸ  ��%�βb�ʸ}g!����g3n       `�-�T��l��i��Y*��u�nC0�G,�^m�,��['K�����e����'�  �01�ncu�΋M��}r���~|�ʊw
        ��Õ�B8�L�݂~3YgY�9/K�w 5�[�����)��K1]���P�w���s��!Ί�  �X�Vj/K�S0&���Oj���y[��        0f�^��])�>���n�f
[v*��� �ŒR{IV�:00By��L{u[e�>�74�'��\1n  ��b�ج+��ce����       OՏ�m���y��/�[��~�]��$�DX�VlT��Ɗ�{�l�i��]�.�N �U&YZ�+EY*d1�_�X�!֒d��K�RkA�Y�V�T!�n��|�%��¿x        ����*+�w�t��}»�$v�5Y��.��eiu��ZX�R8)�^���`�;�D�񼛶��$���,�R\��������7�MV�$)d
Yi��L!d�����ߏ��81)*u�_4�%�\A�U���R�p         I:����U�HP�q�l�Pުl�IǷ  I����Yf��0�������FC�����/��C� F���c��ו��a��%)+����A|I!+Ka(~��ϒRg�a;��?�>%\Ÿ        <ؙ�߰�jf�y�`�Lٖ]
ۼK ���B��$E���l�)�����w{�ܯ�pB�]�n����bWVt�>f��T,J1������4~�P(��8��v��}��d��q;        x(w�\�с��OY	J�{�`�XRj/Jy[��'�>� Ɖ�RwE�m�M0LR(�KIz�w�����߰eiW�����- ���b.+��ؕb����)��ʫ�ޏ��!��81)*u�1 �?�=E/f�        չ���t��.�N�f˔m�;��aEg�j��=��M����������0�Ż��3[��^�eEW��U�F�Ri��;���B�m�����v        �F�VʧnMT�%�)pP�Ti�n��]���K���]`#B�q���=��n���"I�w��)�Ի��2Y�Vj-(��*�������LJ�,o)u���5��Y�Fm�˼%��:s�ւR���v�P~?�v        �f�U�Z;�\��;bw�=�nC��	`�X���Re���;��w��q���h๕�;K�v� �Ê���8�ɿ��
��ciu�^tVG�ݦ,v���ٻ�8I�����s���꽧g�F�4ha&`�5��1X2��%�^/�A�B�˵lc_0\r�k�Z�I,1�#;�/c�q�H,�@ �4�]�{-O=�������MU������j��=�|�ݵ�|�_�%39�$7��@a���ٹ}�kܾ1@�Ǫs~\w���u        '�;Bc���:66�,9�(v��Iy*�R��(�4w C���B�Xl&�l�����C�	����>I;b� 0 �6���Wh,n<9b�n�l��n��K���7��K
�5Y�JƓQ�����P����X��x�`��Oչ�[%�!        x���vu����?����B���\���ar��B�*�v�4 ��앱#5�w�{m� Ⲑ)4W:e�֊dy�H[�岬)K�5�kG:o��\���R�g�S���xs���8&���܁��        ������%op�[bGA<��_UY֌ N��BkM����݈�@��������cH^p7sW��  ˚��5��Y�.���B�����벼-�r'fcZ;�q8s�Gjs�wPn        ]u�u�����7ǎ��,��{{cI� 0 k��>/K�D7������CHR;���}��>S��R� ���M��R��ʴ�!`���y*k7di]��S�M�yɹ�!1 ,d�t]��ܙD�m����U�;        ؤ���o~�'��I���qQȎMCvI�c00,K��)�[�s���>���cbx\.��� �e-�֚ڱ���X�잧?�uI�ExR�KJrIA/ȷ��w�!�i�4�	1���U���9        �&W�����_&�7ǎ��L��)o7�G&䊣���,d��Zgx!�-�BxY���cx<&�&v �gYK�zU��H�}��\�5e�U�zU�����Bkuc�w���f�y7�ƒ�y��2�v����*        lΪ��Er;	��
�e���,d�� �j,(4W֫�ہ���=�����c�Ȃ��7�?�%}O� zǲ�Sr�ؾmLyO�7
�G:%�Ʋ,���x[�!d&ˎ/�/m���g�!�
��¡��c�         [�-��Չ��A�;
D�*�W�+��{f
�5�k�v]t= �к"z�����h@�8E!Wh,)4jLt��,�e����S�7^�[������#'�7����!���zYx��x�        ����jCo�����d���t]Nt��B��|}^�����c�}y�.v�ǲ����kb� �M���e�u�dO����\R����y_�j˱�ɲ�,kq�
6��Y�L?�J�(        ��*��e��\���Q0`\"?2!W����3Y��<cy�0 R�Vm�6�Q�6�v�
�g\���ԕ$����;,KZ+S��u�X��%E�o����=�/�B{�ʲ�6�t�K�x�2{�v        00���f��g����` ���Ȥ\�;	��c�vS��F�����K����{��n�mۍ\.����r�֪,k�N�M+Hy�)_�������^���h)���Lʳ��4O90���ua��7�r�v        08n���k+?0��os
��&�5))u��I1v" C���� NJ���(�e�]-����
麬�.�� "Y���鸇���w�<|�4�oh�dy&m)ow
��m[��OT'/�N�\ǫw        0xn����?x͢j����q0��T�^����	�� �e�p�$Y�_s�k���u݇7v OQȕ7��<��8q.�(�'��DrGO}�t�΂,�Ǌ��g�.��-�\r�V���
��       �@�`�Gj�p�9Qr�r��\i��; I�e��b{;v C+inӶ�{�~�c��*��x�����s xj��Ph�����\�t���+�'�sr�wJ�.�C��)�Ǖ�s��Evn����'�G|���Q^�       ��pƵ�����^;�@2"_�+�b'�w&k7�:�v ]�#�X��=���w!Ʀ���;����BsE�5c'z�6ަ);6����\��Qxw�?�N���D�x����l����ce�����c'�H���q�z�Qn        ��۷�\���T�73�i����y0��B�%��|iL�Xր�@�mf
�,��X� �!/�D�]fW�|
.�5�+L��+�o\z�����ym\?�[*i�,         '��*��/�\F��Kᅱ�`��BsYj�ɕ�䋣��l 6
i]֮���&{I���N>��m�4/)���	0Sh��ڍ�I  xB&�7cӯ��-?ǃ        j;���������];���+����
��a ��SYڐeM1j@o�z��i�Q���s�7|<嶽Z�ہ�`!S^�Qn �?|�q%�v        �,���ms�e���Y0lL�55�k�
��ء �(3YZW�^U��dYC���^��Vz~����n�폝������^�B;v  ���Rh�^�p믯�N        �-+����v��2�;���֪���΀ô.Y��
�c����\���Z����\��"ƾRp7'�ձS x"��ZSh,I�E `����r�U����I         �m�3�Zu��J�{bg���S�֊�#�닲v��;[��u��
���]}- �{I�m]�Mm�>|���s x�7���;	  '���륇?]9;	        @/�\������bg�&�r���GR����,Ȳ�B�IG�@1�j�i�*��i3�}���3 xl����Wy� 
f�J
���        ���C��f^(���;6�Ж�k
�jg�tkU���,v2`� k7K���� 0x���������}��n�+bg �ݬ�P��$�cG �I��7���U?�����        �/˷]����4;6����u�FM����E�t]��ɀ�cA�֕����-k��G 2����3z�}�����c� �H���9*�'O �!`�&I���*ߊ�        �ߪ��r��+D�=gRޒ�V�:�Ʋ�ݠ�<�B��|��|�BkecR;�, C�����ܓ4y��b� �2�ƒ,]� �br*�_5���         �Ń��\�_irK��`�\�5��ޛޱ�Y���
���mb}A�Z�B;v2 xJ�����3z�]�];���7�� ��gr�W�n{ם��         Ķpk��\-i5vlQ����ޏ(4��uY����؜L��
�����7�d�dy�p p�,���cW?��^pw��3 �N^�Iy;
  '�䖼W,��cg        G�n��T|���� � ˚�֪B��|�����Bs�)��1d�d�F�}��:�k�t�)� 6+�������w�����tv� $��
���[C ��ox_z�����;	        ����]��·kej��<�I�-k���:��^Sh�vJ�y[��1P,Ȳ�Bk��	퍍B;�L `�0����~�~n�h.	���? ��M��x� �IR��#����Q         ���������()��x|A�SY�>���r��9M
_z�L��e�-�����N �.��vQ'�K��;��u��(� ����
?z��{>;
        ����;��N�OJ.�����ɲ�,]Sh,mL{?�|�ڙ���˲T2~��Y�e�B���XV���|�pg:{kU�5)��g�su��};h��k��R��]w�:,iG���uYk5v  N�����:���I         ���7�����������%�ߓ�ˑg�">3Y�:M��c�98 N�/�;�_��^�޳eǗw<G�ہ((� �����Sn        8y�C7|`��JY
�;��<=6l��I��|���Q��}D��3)Y�%�7���F��)� ����6w�ݛ�<���VZ��t=v  N��Wjs�ߎ�        `XU�*��}e�~&v���Sp�sY���cS������w� ?hl��r�m�n�r=�� �.��"I�ۏ���%��x{[Sh�����1  89��z�P���1         �]u�������_���L�V�8��7�䑅��;��ƬSX�Й����)�@lf�y����k��=�ڛK�n�&i<���V�˲v#v  N�s�?X8t��b�         �<��^��?t�;	��8/�mߝ�F^�s�{���5��If���q9<|���q�C�b ����ON��/��z�(ܫI�{(��a
�eY֌ ��✿y���o�n�        `qV�W���Q?!���Nl*�Q����y�O<���{��9u��������ٶ����;����݉��w���Wظ��p�=<|�	� ��%��z�����FQ
�y�WFl9�� ��T8T��M��o@         ��J�m��]�ڜ\xy�8 $)t�����S�Q �/����(�m�L���/�Մ�
�v ��1�gj�u�uy�,         ��=s?��M]#�/��  ���-<�/��c�����������/�Մ�,kĎ �I�W.�ktK%��        `����������;cg  ��3ӳ��O�'���_$���}�-$4Wdm�� �!c�+iA�y�J=v        ��b�����&���Y   0�̞vƵ��6}/���K��'���֪�M/ 0\L���ܫVo�,��        ����<�
�����   `�9+���K{�M��A/����VZk�t=v  N��#Iq���\�۱�         lU˷]��D�j3-��  �f�z�E_�O���s���{[EH�e�Z�  �$��br����'v        ��n~�/%*]-9�:   ��ɞ��=�B߇    IDATZp�w��K���V�uYk5v  N�o8�k������I         �1�{�Fο�L��Y   0�Bxv���k��ɾ���[���� ��\�Ľya�         �T=t�ϼӏK�cg  ��qn���9��}-����~�lv��
͕�1  8I.x��U?y��N        �Ƕ0w��K~1v   +Ϯ�ua/w�_����Q��69��
�%I;
  '�����^���c         ����-��_�s   `�x����{���v$�K%M�k?`S�F�=�N ��qɯV���1         pb�s�w��ߏ�   ��,<����������~�lj�7%�c' �$��W���)         pr������q�   ��^�޷����q/`s2S�X�B;	  '��iu��O�N        �������?;	   ��^.߿������I�沔��c  pRL�s�4�f�Y�,         x�n��#]#�/Ď  �Ȝ�{Ƌ��h���K������ْN��^�f�+��;  '�����+���V�,         85�V�r]-s���  ������3{�x_
�!qLoNAH�e�z�  ����
�+ks���Y         ��?]9����&�@�,   ��y=�Wk���nο�� ��eMYk5v  N�|�/�~�߉         ݵt��L�6�r�,   �äg�j��eF�x
,o+4z 2��������Q         ��s7}�%��Ԋ�   �gf�j��������.��>�fcA��$)�N �	3S�9���*;         z�z����>�QIy�,   �3��z�t��{å�F{�����ƒd�� \��ma��m��         �?��Ŝ~>v   ��3;K�VJ�X����酽��lBcE���1  8I�����o�         �ڡǜ���9   �GN�m��i�X��w�����LB�.��c  pRL���s�_��         q�U��s�?��  ��)h��^����w�DY��Z��c  p������\�         �ka��w�ܡ�9   �y�E�X���=�~p�L��r`���)4�b�  �$��T�<�F�Y�$         ����r�]+�;
   z��.�ź=-��\����MÂB}QR�� �f�����?ڎ�         ���*����$���Y   �k�^��ӂ��{^/�6S�X�,� �fr��x�­��;         ��m���_m�cg  @��׋e{Zp�܁'ZkR�Ǝ �	3iQ�p�§��_H        �1-z�7gWI~%v   �s;'_����^��ܝ�����agYS��ǎ ��s��8���m7�;
         ���M_rNo6S;v   �F�.���=+�Ͼ��S2]Ы��ag!Shp�2 `��N���*;         ��¡�'��C���  ���ޝ��5��౅�¥�\����)4�%��A  8aA�_Z8t���        ��2���%���s   ����s��f�
�ץ�Zv��"�} 0L��,����S         `8U�*���b�   @w9�s��f�
�f܁�bi]�nĎ ��3�gչ�&v         �����n��;   ������=+�Kzn����m��j�  �03�w�M�Ar;         ��-���D���?Ď  ������fO
�����˒.����в��X�D? 0,���vz�}wT���         `sx�J=)��4��bg  ���rgH��v��\쨵f�^*�bm �ęF
N��TNLEo*%R)��T𦂗
^*�Οi�/)�Zr�F�G��$�'/���{��̤,HfR;�\�N����u�L;Hypj�R����)R�w�� �t�C��ի���j�$         �\����ó���j��wҶ�y  ��9�R�4Rt*x�b���
NŤ�Q.8�TH���JI�[W.:I��:�.(礒7���V�����?Ƕ�IfA���̔�S��������_���ܔf�V�Ҷ�Ly0�B/�]@|N���:�6�owkɞ�]�?C��������i�`-H�E�hb�N��hQשSfOL�S��n4�'���~����;p%��~�3�G��c�O�Y���ʜZ���;��V����S#uj�N��R< l�·���t_�          ؜j��t玫��z��!9+�� ��ђ�h�i�$��x�}���q~��6:|N�%��	�}jN������:�a�y���mS�mZO�9���iP��c�k�M�4���,P��p�!�����%����$��Ƌ���i�d/�L%�XQ��(��M�O�a���jtt�?�m8Z�7�G���~����=���_������:����z*�gN��z۩�9��N9� 0t����޸p�/��        ��m������Ɵ0���d'� D֙�>1�59�4Y���*{M���JN�#N�E�dOos��/���0^���=}ty�#�TϜV����i���2��Ak-i���
��)�#��t���vk���M�lλ���fF��FL�#��d�4U
�*��KOm��fs�S�����<�ef��\c!(<�� [��z[Zo{���ն�J�S~�  �ɹ�g8;         ���C7���+*���M��  ��xM�M�z͌z͔�fƼ����G�Fz6iR�����i�(i����N�-�bӴ�0�4�VZ��f�r�s9�smփ0 �����zRp7�^���c�h�)�fF�fFL�#A����H�x�;�~:Z�O�D�b�	��h�=���d�<�T��B�_�ȜVS��TZj:-�N�-���w ����v����        ���z{��ۯ��/~,v �j
I�m�^�ƼfǼvN$�);m��KO4i��נ��4]���N�q��{8�Z۩V�Ճ�"�b#�J�TO�d�����x���\����?������^�O�K��m����r��i�l*x����^�{
�}�rt�������G��K��>kG���r�i��Tky���
 ��o����T�         [Pu�n_��,�^; lF��D��mw�1�h�������E�Ĵ�Y��O���Ms�jݴ�4��X�U����@a'&�;���u����'/�
�}���rA�1�}̖M�GM�%���j�s*
�[�Ϗ+��e������z����5�9mz-6��m�S�0���ra        �8n�.����|���R�$v V�5;�hǄ׮�D�'�vOx��b'à*%��&��&�:��;�>��Ҕ�릅u��Z���\���v��)�8�s�����^p��_"=��R`�J����c�Sd�9f�14U�N'&I%I�]�?�}<˴m<�YY�<oK��I+-�j�k�鵰�9ߦ� O���+���;*��Y         ��-�Ż�g�|�������;v t#�D;'��L�g����f�hp�;���4]v�`֩S~/�LZiI��M�ׂ�W�փ��߷0��s��ߏ��C�fҿ���,傴k,�=�]c���M�GF���)˲cy���n��d&��NM�j�k��5�p���8&�$���*w��         ���+�ɇ��4; ��B�ݓ^���6�h���(�=�ܤj]z`%�C���+�փ�,�޷ SV�?8�/~�ݍ�~����朮�����������=�g,h����؈���#���v[!t��-���^Ն��F��;���L����?t��          �������͒����`�s�kf�Sh?s���f�vN8&�c(���+A�=����Z�z+�������ڧ��n�U��"�s^��;7�J��g<h�x��ƃN��*��pI�DI�hdd��uGK�c�Of��3���B��H��p��uϔw [�%J~�r;         U�`��WU��B���Y ��F��N�Jt�L��3�t*rx6�ɒt��wx�-/7��WL�Y���r����,���)3gI�J����\���#+��uq��P�N�V�Lf�3֙�~���;
������n��e�L�R���z����z����a ��z����1         �'3{��~�Y���9 ���J��Nt�t���%:m����ڂI�u�wV�\���J��Z&3���go\������X��ܗ&
�x�����N��;t�dgB{����B��B��r�,I23��m���vO����r��u�ֽ\K��@1 C�9�¡�$UbG         �T�2{��߻����� �S5>�謙�Ξ-����1����vN8�H���:��V.ݿd��R�o/�:��)���I�D���Z��w���GK��i�x��A{'r��O�9�R��R�$�Sx��\��vM����Vm��������z��z�����'����          C�R	��T^����H���q �D�ݓ���^�y��N�trtځ�2�Hlw�`{ARA�FT�K�Z
�9��K��mI�`��խ��Zp���{����\gN�:s2hz�p*�sǦ����J��,�d��S�.NS�����zp��;k�Zw�T�����;*��A         ����m�����5r���� ��y�u�T�sg:oG�Sh�
�d��v�K;ǽ���K*��(�Šo-�1�Z3��x\��Z��w����蟉�錉���r�3�Sh��
�Si�3fR=�������}k�龕D�m����L�r����*��          OEm���WV��_K��� &G�=��ق��HT.��mvT��z����RC�����L��r�2Ὧ��-�;�Îzg�h:{�3����\3ent@lG�ccc23�i����ΚI�¬�Z��۫N��$:\�<T�;3���ks         8�*�8{��~�Y�ǒ��y l-�{�Nt�lA�v�s��$0hfF��Q�g�)�3�}T_���f-��˹-&���3�޵����$��Cw9��n�����w"�9ӝ)�ǂ����!(MS�Z-�ig���뉾�����Di;!���\�C~'v         �[���=��;��o��uֶ��ߑ��]��;R@�-6�{�����V��<P��&᫵O���n��ź��]�}x]�h���zfʦ�3]�-�ɠ�q�����,S��R��R;�u��u���}ˉVR�^����s����         ���+�Q
o����39���ق�����{%�z�M)��+N�.����L��B�X���|����V��w�x�����^�@��$��s�3��1�}�H�،�s*�*����P��j�tֶT��S-4��[�o%�R�g� N�������b'         ��:��Ϯ��cg0�v�w
��L�k�ǎ�
^:w�t�LARAk�ӽ�\�Vs�W��J۱#!�Mz^A��)�֢�q퇾�;�ѭ�6��A��:g:���\�.+������Z���4U�!ݿ��+^G�<a�T��LzQm��;	         �+�W�k[!�>/i_�, �϶��.�U�3v�s�����I_��to5��j���'�Y{`������ӵ	����2���Hb:g:輙\�M�gJ;��x�U.�U.�ef�JS�6�ҳ[--6�o,'��r�E&�81�骥�)�        `s[>�k���+����uNӱ� |�&�z�΂�������i *��&��&z�y��e�S�{!ӷ3��Lw<��������-�ӝ��}�Lٴo[��3�J�8�9���hdd�X�}�LK�KS��ҽˉ�]J���N
` �k&.����7�;
         ����]��������rֵ.��c�X��v���=�����q �ɒ��Ӝ.=��<���1}m>�����$��G%���tq�{�k[|���Ѡ�fs�?�k�X���� ����Sm�����Z��M�,%�{��F;)�a��w9t��b         �����|jە7��7�^�, �x)Ѿ�]����g(���K�m3��-�O���������S=���,Ď�?Ӎu�8�ݝ�-�8���ɠ}��.��5Y� ��S�TR�T��Ą&'S�6����i�;�^__J�e���!`�rɯ�:���1         ���o��r�,�3v q��};Kz��E���o�:#�Hv�K;ǽ^|vY�M�+�A_[���R[!����y7Xw9�޵�X��Ο	�p6׹ӹFڤ �����驖����z��olLu��St`K1������N         DS�L?5�y��)�*v ��t涂�uZI��*&tf �3]�^p���,����kA_��t�B�|˔��t7V�^�]���^J��3]8��������`08�T.�U.�5�f�[�dWC����(���c��[�F'�Dr<A        ��V�������tq�8 zgz4��w��E͔)�<��Y{�����4/�����m}��V�e����ug�{w��+��]MIŮ�7 F����ؤ���� N\��j6�j4��β�k�����(��
l*&����js�o��         �]�o:?S��N�;��)&^�v���%�=C��pʂ��U�]G2}c��v��&ؚ�j����NW&����ޝR{���#�i߶�g3�3�+��`H%I���q���kj2չ;�Z��t�b��T-�x�=�2��r;         �HG殿w�����B~й�3�تv���%=�D�� í�M�.�YP
��6�;��z��v{Lv�0Սe�Rp���k8���3�3�)�_8��8�� �J��J��&&��O����=���Z�{eLu��y��9?W���A         �AT;t�Ϸ���H��bgp�Ӆ��z��%�=C���T�҅;L�(*����h���>�*����"78w����(�s�r]�=׾m�J	�N ���^�����T�3gzA��{jNwULu�������+��         dչ�q���[cgpbvNt�ޒ��'���l!�3훕���|ZQ_Y�ݿ��VCTv6ݍe�Rp�޶����I�;�)�_�=�h�R;���P(hrrR�>�ҳ�4���\_�t߲����2�o��@���c'         ����9���������y�oGQ�sfIg1� T.H�����=%��Gt��\w���r*�;����2])���m��o�>��.ޞi�De ��S�\V�\��d��v6T]m��U���
jd�x$�U�~X�ʀ?S         �?�n���b��d�Ď�a�D�>���Q��Ȁ ���3�.;���fI��P�;ʴ��J8��9W��:])���3��M+J϶��������qt�����v�4��Ӛ��f���h��ѱ@l&-&ő��o}�J�,         �0Y�������q�}N�d�<�V�w����-��yz� p¦��K�I��s=�V��| ӗ�j���ю1��ܝ¬)�#M�s�r=}G�}�r%<��S���ؘ���45���=����'��R""0�%���[�}O�(         �0Z<t�?︪�#�'$%�� [�s�;F�³�:c�A� p�N�0���D߿oT�\��|�������Y�\f68wsn[��������_�#�hap���fP*�T*�41���ن��-}y���jAi;�u���v������         ����[g�Wnt
�*J��%{Jz�9EM��Z ��t�t�LQͧ�Յ���;�R��=G�~����:]9q쒫��szZ7�:A:�ǝ�o����8}Ҿ��A] �3�{�J%MO���i��[Kr���Z9/>��r��U�;         �4�����|�dϊ��̦ˉ^t��^�̲.�U�H�~	 �Z�K{&�^xV�ѿ9<��Ω�L�da�_�,m����^:���]����n��$ڒ:����Ço��L����>� ��S�\V�\��TK�����2�ӑ�(b7    IDAT�M^� �f���6�࿎�         �L&z�꨻X����l6{&�z�9%]�+M ��9����?U��sz�G�ݮ#k��Y�m
�岬+�џ`��t�]y�u݇�Y�3��֣9g_��>�B�?�/o;|��~�7�"I_�ž ��e�����]h럎��:/O�n0�[��?��+Gbg         6����3���퉝�Ι-��t��& '"H�����_��u9M����o�<=���?&���܍�6ʺ2�]Ҷ.�sԚ��l�;������}����9�� S�P��Ԕ�5�k߮��Gݷ�cG���{^wx�r;         ���ʷw��r�>#���y�a�Ӿ�E}�9#:m� of��t��W.|�J�Q��v\��/Us��Ph�ukc'�t�9��/~��Ic]���������.���O��s��ζ �S�$�&&&t������Ѓ�}�׽��B�p�p19����          �ّ�>����,�p�,�0���{��޳��6� D D�糶p��J�_m��#�I{��-K߮�}�����-\\��橬ѕ��I�S��-'�*飇o~�_���T*%I/;�} =����ؘ����-Yj�2}�Z��� 3�[���9v         `+X8t���^Uy��m�� ��{�Kv���J�.3� �	_��˒~[�oo�o?_y���?���>Ս�Q�<�?{T��z*�����b;�=|�;�;�r�$MMM�H��S� ��9��e��{F��hLo~F�g�̔��x��w�і���w���]-=XT�# }�"��51AA��c<)-�x�j��Z�C��kNr���p\8��hc�����{Q��F���f����D��ݬ�޹���>V��>����6�?���K�yC�      ��L�����\}�t��fU�	ƫ�6/8fH�`~X�q�ƣfr���x��'>�_^���jp�?Gc蛳��w�ι�ޅ�9E�g`�ޕ">q�ͯ�XDʳ��n��Mɍ��)�?ix8�Y�3N�{��Os|cK3ڳ��s��ݻw����.�      �/����j�pw#��"V��u1Ш�����kc�R;��SUչ�^�o[�������w_yjx:�w�c�7���[�Sn�+��_�<�����>�r{DDJ��r= �744�"~󨱸�v�w�Fw���i[s0^��co�(      �{?Һ/��#���@iͪ���?z�X<��!�v�y*�t�\�xd�{sh�Ս�%����]3\5缀}�w�}^����������v���} >њ��G��mo�kpp��BA�rv��[����N|��ftJ�2rj^��k��t      X��yΛ_�I�,�JH)ű�obc;��uɒ%{]~�廻vb�U������w����ψ���Fg�OW?�鿸k.c�ܐ���]��iG��%�������W�z��<;������8p���{ٮ8~����{r|{�sz��;�u��      P�߱��z^��ȝ?*���J)�� �>t(�)�,$K|��3#�S];���������^����ij�k�ԮK��{����f5����;c�`��"����6����7�jr��>�n���>c�~����q���?	Ew����<#�16�N      <b������zr��9��@o�8b��8簁�k̾Y����:��+�������FīW^t�Սm;.�w�6ڻ����9���|�T4n�����}�Vg��M�o�i }444�����Ll��q?��(�T}'�zI���׿�      ��h�:��j]��_H�Jǁ^8t��8����w��v��,��[���3&�v��#���j�g�-{~~x���z漻;]��GG�7K� ��v��߿������nWtg�i[c0=����Z:
      �g{�N�Լ;>�)��e�%�8爡8dE�t ��]UվW\q�d� 31ۂ� @��OZ�0����K'�nH�\U�)�     @�m�p�Q�WGD.��j�h3~���x���� �K���<�t��Rp��RJ1::��<.>�O?���S��j���/      xb�o���ݥs�l�6⷏�?8s4��G�`��w��yUp�{�;�,���K)Œ�8��eq�U��;��]"rT�8=_[:      0}g�k#�(�f�Q�8u�p\���8��fT�t" 
���fj^ݶ�����"�S�s P^�ݎ{x(��G��֤'���釻w�:u���>Q:      03�?�m�슝_J��T:<�#��s��eå� P�F�u��}�t��o�o�U:  ��h4��������c��\:<��᪙�Sn     ��駛�xJ�EN;Jg��r�����x���� <Z�ݞW��Vp?�t  �e`` �<pY\x�p<��v,Pt�~RJ����R�      ��MlZ�O��ה��j�p�۱�q�)#q���V	�O�{��jGę�s POCCCq��q٩����10o�p,t95޻eӆ���      ��䦷�YD���s@DD�������g��S�o��@�=;�J���yS�FDxq
 �)��#q�Q���8|y�t$��+�זN      tϒ��U9������v�>C�O�s�fc��(g�o���!�k��SJ�� ��PUU��x��	K�G�X>�KGbQ���4����y���I      ����'Z;���H������=ֈO�?ˇ���v�����k��s��*�����l�q��ť���������1��4�S��[[w��      t߃�����^^-N_5S<��x�c�z� 3WUռ�bϋG�6nܸ��hLFD�t 槜s������N�][���y�ͫؼ���9      ��Z��7�%E�M�s���P<눡ў`n<����:���k��޼x����g�r; s�R�V�������|(��ĂU}@�      ����7�T�^:�^c����x�����ew�u�ɥCL�|)�ϛ�� �[�шc��4.;u8�vP'�ŝ�y#���KJ�       �%��qa��;���p6R<��x�cq�r� ��٥LǼ����誑�8��eq�	�8x�m�tC��48���?��V:	      �?��[?�"Ώ�.���������*�N�B�R:�t���-�mo{�^�����<)�0�LMM���=>��"�]:�T����ۆ��t      ��}���WvR�/K�`~Z:\�o5���(�,��}```�ڵkw���xj_xṽ� �_�f3N\�4^q�P��o��OQCջ��     `q���Q�u��?�0�:cL����9�NMM�Y:����g� ��0>:�9vi�wl#��N����41W�N      �71��T:����f\t�x����jZ�@t:��w�k_pO)�S: �GUUq��c���G��6wW����L���v��      ��-�]�j��9��Q���R��j8^y�H���> ���ͮuo��ۿ�������s�M|kW��p�o��:)�nټ���I      �zY��7��r�戬�̣�5ֈ�3-�� �쬪j�W\�p� ���w�F���3 �x����F����'�z�4�՟*�      {2�i��s��J�>U���W�1��@iC�v���!O�NG����qΑ�q�Ƀ��X.�Z�>6�y���)      ���<#�̩�T�����f\v�x<�����@������Z�SJ���`�H)�+���S��7V����^ʑ�i���i      ౵Z��=𒈸�t�hT)�:t$.;}4��l�>rε�h���y�M7�k׮{��X��}pG�ݿ�os�ZLr�]Q�3y���-�      ��~�[��c꣑r�t�g���x��C�lD� �Zڱm۶�VkG� {R����w�>;������ǅ���9�T��/&��F�      ��-w��9�?)���jV�ܣG����������SK�x,����}�= 4��8������8`�tz����7�N      �?�w�K�js���A˚�3��ăJG�'�R�mW������_ ��}��E���%�Y��更헔N      �W)�޵��qW�$t_U�8�������X>�9 ��P�e䵼��p�+;���Q�> ���'w�m��#�Y�[,��cg������JG      淽^��b�ԧ"�P�,tǊ�F��ؑ8h�� �KJi�֭[W�Z�]����Z�U���3��� ��<i�P����8q�#5�)�      �0q���w��s��0�<}L��y)�<�dɒ�K�ؓZ�YSJ�]y Odh��9f<~���(��9�Շ&6oxO�      �����6�H�J�`�F�������@�t ��N�S��v-�qv�  0)�8j��x��q�J��磜�t��/-�      Xxv��uI��Q����{��9G���������v��w��˚��DD�  B�9�|�����MŮv�4LK��1�|�ĭ�?_:
      �0�|��<-:��L�Kg�6�8���8m�W���lݶm��V�5U:�/���F�qV(������U�q���q�x�-cOR\��      �����~6��U:Ol�%�x��c�� ,DK���O*�Wծ�^U�3Jg �^�{�`����8kU��+T�%Շ'6���K�       ��Mޞ��\:{V�g���N�����`�:�t�_U��{���3 @�4�xƑK�%�Ÿ���N���qq�      ��{�΋s��K��і7⢓G����m`�cw�V��n�i("N-� z�}����ơ+�\9v�Ըprs�祣       ��֏�}��r�ݥ�������>OZ�( z.�d���ٱcǩ1\: ���P3^|�x���j���T]3�i�?��      ,>�m^����ͥs,v)�8��xɉ#1:��| �����#J��e�*���	  襪J���F�'����˩n���zW�      ��5���o�)�Q:�b56XŅ'��3���{ ��u��Vpz� P�ꕃ���b��Zݚ����t      `�Kyw#]�#�]:�bs�ʁxՙcq�
���8UUU�wm��9�O-� J�ₓ���C�s�^�r�j�t��>��Y�(       [ommiF��i�t�� �g����4�ֶ�x�k���Q:�#�,YrLD\U: ��R��Wē�������.�h�K՛�ln�M�       �x�w�h��sS�KgY���F����� �׹����~���Q��Q��? ��f��x��c�zy�n�L��ؼ��c       ����cC����9�5+�Ug�������"��C<�6w�sm�R �Ƈ��ऱ8{M�>7�"G����)��      �kZ�Nj\Q�_:�B�R�3W�'��蠽� ��RJ��rצ/W�� ���J���F��c�Y:�B�:UU]6q۵?.�      �L�v�#w.����`l��4�>�� �Gg���Zܫ�������I� Pg?����O�uJG��rT���ZW:      �t����{"w�S��فK�q���1>T�}� PG��m۶��jm/�w쪪j����Z:҈��:'�(e��9�29W��      0]c��՗K瘯�;`0.:eD� ����%K�("�&����Kg ���٨�9ǌ�o9�Z��e>�~�h�8ni�*�      `�ni�F.�����2�TU�s��3��� 0M�XZ^��{��i�3 �|r��x��#16���"��ۛ�S:      �Lm����JU���9�с*.<i4N}R�t �WrεXZ^�w�7�t:��E�`�, 0�<�������w[�t�zK��Llj]\:      �\����-�鼨t�:�I3�;~$����|��m۶��j��Ҋop�t:��r; �ʲ�*.9u,��o�t��J�w�����1       �*w�9��K稫��KNUn��[�lٲ�J�(^p�9?�t �Ϛ��{�H<���f��;�Q]t�'Z�JG      ���ͭ�Gn�,��]:K����G����F�F �o�N�x����<�tf� ���z(�?q$��j�ȍ�ډ[��t      �n��c��"5�Z:G]�T�ғ��7KG���ˋ�#�� `�8t��x��c��xn������7���1       �mr��?�\�Y:Gi{�5�姍���#�.*�������_��  ��*.9e4�ާQ:J19b"�͋#R.�      ��R�f��iK�$���@\v�h,�s �c��w,+�h�=�T�� �@��>e4�Z3��G���z��m���t      �^����W�Z[:G���♇��yǏ�@c~# �W5��Ӌ(9<��Ԓ�`!K)�3�7�����>W�_Nln}�t      �^۲i��"US:G�4�x�q#����� �BW��]����� ���`\x�h�.��{��3\��J�       �j{�:"�W:G��T�ғG��}��� �bpf��Śn7�t�Ю]����R `1ypG'n��ñ�v�(=�#�J��Y���|�,       ���3#w>�R,���+G�Gb�H�}� �h�l۶m{�Z�N������w�>%���o�Wqɩ��f����R�Rn      ��ͭ�T��t�^8xE3.=mT� �k���������真Zj6 ,VC�/9q$N8p�t���Q}rb��w��      P�����gJ����N��f* ��]��Yp6 ,ZU�xޓ�㙇���9�h7_�r�,       ŴZ�Nj^�#��t��Jq�!��c��Q)�@	)�b]ow X���f0~���h��5R�?M~����      P��6]����xM�sѬ����F��.�7��<T��]��o��v�}O�� ����`;��W��C����\�?w�^^:      @�����ˑ/(�c�F����Gcղy�� ������׼�5��=�ȿ���%� ���e��䔱X12��AN߭v���      P7�H��H?,�c&V�6��S���F=��I%����i�� {�|���N��+���LW������Vߟ      ���ͭ�Gn\9M��2�V4����b�|[� \UU��[bhD�� �mx����8��7P:�4T�ۼ�3�S       ����?��]�s<�����8��f ,*E������sNqJ�� O�Q����F�����8җ&ƏY_:      @�M���7樾\:�c9u�P����hT�t `ϊ,5o�{�ҥK�����= ���+�1�H��ɺ���z87;�{�|o�$       ���/v��|�gS��"r�^�}�������| ���{�{>�я>�ϡ}����� �̜�z0~���EN�i��7N���o��      0_<�i��:�j���c��<�~�!���  ӐR:��3K�O+0 ���n�Yj�FD_��۳�&7o���)       �6�靑�;K爨N�:�)4>Z:	 0=)��/7�{�=�� �C��n���o������
�#�/�H�T      ��+��@\�s<X*A��`���'6�>XU��J�  f�D��������qb?g ��񫯾�����6������o�~R"HjT���ܺ��l      ����[[wU��k��龪�����wFDLMM} ".� ����������>%"F�9 ���ң����C�|-7�̈�[��Q�<q[����L      ��h�m�6��@_���ݩ��[n������zk�yS_s  ��R���o\�ϙ}-�7���� feWJ郿���ںk�9~VD��=]�}�Ow�Q��s�    IDATf      ,|�;��~�ʩ����Y������UU��=] �O���k����Pp�y ����+������s��T��̈�=NѩR��[?�Ɖ��      X<~�w�ɪ��srT�ɻ�~��������n�z{D<�� @w�n�=�|z?� ���O��KkۊX���Շz� ����Mo��g�      ,R[n��)���݄��������,��Z��ko ����[��hD<�_� �Y{�����D���;'Όߏ����G��32����?      ����FzmD|��禔�r�xQ���5��?��5 �RJ��Z�����6hll섈h�k 0;)�]u�UM�íVgbs�9һ���su�ݷ\�p�      ���skk{�/��v���Uu��Mo��h�:����m�>�vk> �3�###G�kX�
�qJg �7�'�'7�y]��-��Su���?׍�       xl��q�sTޝӪ��������Vk*"�ߝ� @/5���5�o��R��P ��=�u�֏����ͭ9��8��+��7��       �ie��&r�׹���Ӊͭkfy񌗰 E�m�y?7�+�@ͥ��{���5��'7oxk��ED��9��4P]���kw�v>       3���kw�@㒜c�,.ϑo�ؼ���ο��+??��� @�,��Vk8"���, `N��d��ۯ}WU�6"ufr]J��|�����      `f&n]����fxY����6�}.�SJ9"n�� @_��sN�ԗ�����S"b�� �Y�oժU���A����?���ў���'��[�1      �����7圾:͏��j��6mxg7fWUuK7� zjٍ7�xX?�����i 0K)�����,�?��7����j��%�iWjƥqKkW�f      0C_�����tq����l��x������n�^�n�SJwu�< �7������ӗ�{J�/ `�r������~�_WU�9���ӟn����n�      `f��p�9U�9MEռl���͹)��s�P7� �/�ԗ��6� [�m�vg/����D�.��S��K����i/�      0s�gě#W��W=�؝�ꒉ���M/榔��� 躅����j朏�� `Nno�Z;zu����3R�pnv.�[�o�j.       3�juR5xqD���/�H���E[6mx_�ƮZ����W� ]qJ�9�zH���E�P��  ��s�����6|(�ꅏ�O�NTo�������\       ff˦7~;R�'�����λ����r���ߎ��z9 ���_��^�y�=�tJ�g  s�shh�~��c��E�~'ru��w���L       fn���1��X��y[6��R<O)�|9 07UU����^H)�� ��߯]����6qǆ�E��)�k&       3�ju&"�ѿ�v�n��������_3�;%"���=��'�a 0K9���r;      @�����V��#���~� f������ӂ��7��H)=��3 �9��o-       ""RJ(� xl)�{=�����눜�h/g  ��R��������       SSS�EĮ�9 �Ǵ������z9����s�� ���=�      @m\s�5��>Q: �ئ��z��i�=�tB/� ��h|�t       �e��@���#�ӂ{�8< 0'_^�n��K�       �_�l6?��9 �=��tw X�<�      @��u��7"��t `�r�'�����o��}"��^� �MUU
�       �R��w� P_G�Z��^޳��Ν;mo����W\��!       `O���; �Wc||��^޳�{JI� jʓ�       ��W\�݈�F� �c�YW�g���: ����6��        �'缹t `�z��w X|�t�       ����z��'�V�5G��l `�>�v�ڝ�C       ��y衇>[K�  ����s���=)�/Y��؈��� ��y�      ��k�Z�RJ/� أ��|�;���=)�眏�Ź ��5�;Jg       ���9o*� س��N�ɹ�8T� j�_֭[���!       `:��; ��q�8�'���z ��ͥ       �t]}��wG�7J�  �h��s�O�Ź �ܤ��      �Wrξ��z�Ig���n�aeD��s�9{h``�ӥC       �)�@=q�7�t��^lp�� ��ck׮�Y:       ��ҥK?�� ������Q�>���v��� ��v       ��/�|wD�Y: �몪�zw�܏��� �5����        �d� �S׻�]/�WU�� 5�s��u�_:       �F����t ��r��.��S���n�	 t�'�      ������#��s  ��RzJ���j�}�ƍ�"by7� �B�      ���w� P?�n��Ʈ�ǻZp���y `��T�       0)%w ��v���yW�9gw ����]�vg�       0��㟎���s  ��RzJ7��v���� ���9�}�       0W�_~���d� ��圏��y]-���lp��i4w��        ݐR�x� ������o��Gu�< �+�[�n��K�       �.�� ꧞����C"b�[� ]qgJ)�       ݰu�֯DĖ�9 �G���|��:�k���1�: 莔�'�      X0Z�V'">Y: �h�F���:�k�N�ӵP @�(�      ���} 5��e�]+�����^���+�]:       tSJ��3  ��s�����Z� 芏�        �v�W~3"~Z: �(����sNqt7� ��+�       X�RJ9"|' �R���ƍWEĒn� tG����<       ��o P;���o_э��Rpo6�O��9 @�|oݺu?,       z!���� �G�J��+���Jy �+<�      ����7��{���9 ���s�J��+���� P#^�      �"��� ���s�� سN���       ��RJ��@��g�{���n� �]���W_}�=�s       @/MMM�}� �����w��]�E�^]� tAJ��3       @����o�� �B�y�ƍ����9�;���� P#^�      �"b	 �Gj4G���n܏�� @���?�       }��� �G����9�s�
� P�z��_��t       臩��ϔ�  <J��)%w ��ϖ        �r�5��?*� �ws�Ϲ�ލ @w��      Xl|W �Q���j�#b�\C  ݑR��5       ߕ@}�sNs9`N�e˖͹� t�ĕW^���!       ��:���; ���u�]w�\�S���n�y�< �5�M)��!       ��֬Y��Z: ��fsN�9�s�
� P�-        �����oG��,� ���v��TpO))�@}(�      �(�}g 51׎�\�G��z �kvo۶��C       @	)�ϔ�  �B��s t͗Z����!       ������ED�t  ""��o�ᆕ��\� ݑs�$:       ��ڵk�(� ����o�ᆑ�^<�{�ݶ� j���ϖ�        %Y �QE��s�xVRJG��Z �����>W:       �d9 �G�y�]�Y�c�z ��~p��W�S:       ���tlp���t:���
� P^�       W]u�"�ǥs  UU6�k�0w�C���5       �w�+  ��9�� �U����9       ��%q PG���Y������+f; 莔���۷�t       ��ϗ  DD�A7�p��l.�U�}``��v ��n�ZS�C       @l۶�K�{t (/����fs�
�)%w ����Jg       ��h�Z�#⛥s  ��Ϫ��j� ݕRRp      �G�]: �@_�9gw ��      ��RJ_,� ��t:�+�϶M t��m۶}�t       ��N�cY �@_7�G��; ���V��)       �䡇�JD�.� �]�|���n�iiD�;�a @��=q       ���j툈��� ĪV�5<Ӌf\p߱c��� P_,        �(�di �W-[��_4���Й^ t_�Y�       ��[��:��a3�f����[� @�=x�UW}�t       �)K� �:�Κ�^3�{Ji�L� ���)�\:       �ђ%K�;J�  b����#b�,� �˫�       �1\~��#�k�s �b�RZ3�k�`~�*5       x|�/  ���^3������ �F�a�;       <����q PX�7��t�M�DĒ� �j˺u�~X:       �Y�ӱ< ��{�ƍ3�Ϩ�k׮53� t]���       �V�^���x�t X쪪Z=����� t_J�K�3       @ݝ����Z� ��UU�fF��ɇs·�( �u9篔�        �����N��f&��Q�=�d�; �R�j�       0TUe�; �7���
��f�� �kǶm۾[:       ��v�9 (,��f&�Wp����Vk�t       �:��W#"�� �Y�y�L>?ӂ��3�< �]^�       �t�5�<w�� �Y�6�_��{GĒ� �(���       3��� `��{�ƍ��O��^U՚Y� ���^�       LS��w� PXUU�����~��鬙U ����       3PU���@a3Y�>�{Jiڇ =q�UW]u_�       0�TUe� 6�e��.�GĴ�� =�n       ���:���p� ��M��>�{�yͬ�  ݢ�       3t���#�_J� ��,��f�����i
 ���J  ���Ǯ�>���6g�CR%[�\�
I�6E��.�m��A����.�`A�ݹ�@S&��WзiP�v
[�*�rdQ_4CΜ�za����e�:�����9$�;ba=��     ��r� ������< <z�8:l      ��Lw� ��#_p��7�O<` ��m��g^�       `�� &O�>P�@�R��* ��y6�m�       �hmm���  S������|�@�q� �ƫ�       ��:u꣈��w ���|���|�@��<�? ��Tp      ������; L�A;�*�GĿ~�$ �C����        ���; �Uk��A�w���A�1 �p�����       `�e�O{g ��;���Aܟ�  ���:y���{�       �%g\ :��u�Zp��Cd ��^z饭�!       `��Z�����}�gϞ]��g: ��      �!���+��� ��w�yg��K�ܷ����h�  H�       ���  6���_��K��K)�� Gf:\      ��ad :�a�n���Z�w ���       #s ����3ӂ; tt��u�k       x2�� tt�n�w Xl�����       �	w �� �t� ���      ��|���#�Z� 0a��~� 84
�       ���f���Y� 0a����< p8j�?�       3�� ��Z���k�
� ��0�       �h���N2s�n���7�x㙈8�� �e>�[p      �G(3��@?O�;w��^_سྲ���< ph6�^��^�       �8����� `�677�\q߳�>þ� �����l6�       ���|�����s ���9¾g�}>�[p�~~�;        <n^}�����9 `�����_y�Y ���z       �ǔ;y �d�/��Z��h�  ��?�       S?�  �����=��/3sϿ �Z��4       �s ��C-�g� 8<��\�       ��9 �g�����Z��; �������!       �q�����+��f�#��#� ����l6{�       ��Q)E� ���l6۵Ǿ�/�x≯��{ ��d�W�      �!y��/D���9 `���<yr�!��
�{N� �ǫ�       �p��~�_��kW]� �8����        ��Z��9 �$3��^k���� �!       ��y ��
�{�% �p��5h       p�j��������w-�����É �^�t���!       �1g� :y�ww ����l�Y�       �8�Lw ��wv�Ů��x��  �s�      �C�����{� ��z����	 8<�֟��        ��_|q��� �����ZkF�- ��R��;       4Pk��u �����z뭧"b���  ���       md��; �q|6���;��qܵ .�g       h#3��@'O=�Ԏ�������Í �f{{��3       ����n� 0U�u�w,�g�w �����Ƈ�C       ���{g ����|����� }|0����!       `
�����3 ����^k�q� 8\�VO�      @#?��>����9 `�2s�����ݾ ���d8       4��5">� �h�Q���w�{ �w       h�]= ��cg}ǂ{DXp�>�      �-o[�>��n� :��*�      @C������q�]� �0�
      ������-��Z3"�p�q �{d�C3       4���� �����x�g"�ȡ� �v�������!       `b��@ko����w�������Mx ��y"       [__w_ �lnn>{���)����{� �Z�'�      ���~��W"��9 `�2�q�{
�a� :�LO�      @F� �w X`�       ЇQ: � 3���g��w� Є�;       tPkug }��^kUp�2���       Ї�; tp��ء ��tX      ���@7�/�G� ����       `�J)��  STk=Ђ��d �t��_��       �h{{�W�3 �D��S 8t�        SUkuo }�]p��ff>�. p��2       t�ꫯ^��+�s �}���Qp?}���14� DDD�ի�       �/�t ���ٳg�?��;
�kkkO�� DDd���       ���= ����uG����˓m�  ��)p       �֪� ����^p���; t��       ݹ���qܽ�^kUp��      �/w� �Gf�����/�6�qtH      ��J)�����G�-����~�;       L�w �cς{DXp��6^{�O{�       �)Sp�>J){�-�@{�       ���֖�{ �㎑v� �Yf:       @g��������; LM�u���	 >�8      ��2�f�{� �	ڽ���
� О�;       , #u �����{��d  �}�;        F� �� �H<�       ��> t�{�="�j ��̴�       ���� ����[��gϮG�z�8 0q�8��w        ���Q� 0A'f�����
�yr�� �i����        Dd��; t��3�<u�Ϸ
�����>q `�677�      `d�;| �`kk�V��V�}Gw h��l6��w        bG� ����H5R:    IDAT
�y�O �4O~      ��X]]Up��a���^J�� ��Z�      `A|��_�c� 05;.���h� �Lw       X/���<">� �&3ou�-�@_��        ���: h��j� A�ա       ���@{;�3ӂ; �g�       ��| h,3o�����\� �s(      ��m� �ގ��D�, 0i^k       �E� ���7������� .�       �X��@c
� � �󹧾      `�x; �WkUp�E����P       �ł; ��� `~�ҥ��C        ���h� �Sp���l6{�        n�A� ڻ��~�����X� �Ɂ       ��˗��@{�f�Y��Qp��ώ�� ��q�        ��f��fD\� &&��׏G�(����D�< 0Iz        vt�w  �����7
}� �$9      �b��w  ��������|�� �9      ��Lw� �����Tp��,�      ���*�@c�����8*�@{�       ����@cw�-�@{^g       �ɝ> �ws����|�c ����        ���*�@c7G�KDD�Ղ; 46���      `1�����Xp��v �)�8      ��Lw� ���q�c ���|~�w       �^�8*�@{�#,�@7+++�       ���� ڻc��֪� m]{��7z�        �� ��촗���-a       XP[[[���=� ����       ��=zT� ڻ]p�Lw h�A       ԩS��E�F� 01��7?  m�Z�      `�y;; �u<B� �(�8      �b3^ �Z-�@/�      `�e��} h(3�(�� &'3/��        ����� �����A `rj�
�       ��.�  S��ke6���8�9 L��;       ,��Tp��j��-�G���Y `��      `����n �f�ّ�����;	 L�C0       ,6w� �������0
� �X��R�       ��J)������������ �e���      `����n �a���󣽃 �9      ��� ��Zp���C0       ,6�u ��Z�Lw h�!       �|>w� �mmm���Pp��������!       ������ ��0GK��h�  01Wf���;       ��R�w h,3-�@�       ����w hlǣ%3��-`       Xp���� ���\+�֣�� ��8       ��;u�Ե���; L�Z�� Ж�;       ,w� �P��h�Lw h�R�        ������,�@��      ���� �̵Rk=�; L��/       ,��t� �Z��R�j�  01Wz        �Wku� mYp��2��       ���;  L�Z����) `J�qTp      �%Pku� m-��� e���      `	xK; 4�Vj�G{� �)q�      ��a� �Z+a� �Q�       �@��? �uT� +�8�      ��v hn�d��; 4d�       ���� `b�J��H� 01�       �j�F� ���J�u� �d�_       X�� ��%3�����m�_       X����D��; 4�����       K��z�w ���J�U� �v횂;       ,�R�;~ h��:��Tp���~�i�_       X�8�����
� ����^zi�w       `�֫�3 ��d�P"�� ��n       XG�q� �Z�Rk�� �8�      ���L� ��P2S� �Qp      �%q��%�� �V)�� �x�       ��l6ی�y� 0�9��(�� ��l�        �w� �H��H��#�� ��l�        ܗk� ���C� 0!�       �\��@#��A� �L�^       X.�� ���JD��A `*j�
�       �\��@;���Z���      `�x[; 4�� -9�      �r1f M)�@c�       �\��@;
� ИC/       ,� Д�; 4��       K$3��@;
� И�;       ,w hG� Z�T7       ,cv �NQp���qTp      �%Rku� �%"J� 0!��      �%�m� Д�; �TJQp      ��� ���w
 ��q=�       ��]? �S���R�C/       ,� �Hf�c�  0�V�^       X.����Z�h� ��       �%3��@;��%�       �\�qTp�v�w hK�       �Hf^� &d�� ���;       pp�Vw� Ўw hI�       �K)�]? �c� ZZ]]u�      �%2���� `B,�@Kׯ_w�      �%2�1; h��Z-�@Ckkk�       �Dj������K�Ղ; 42��C/       ,��|�m� �N-��� �lmm)�      ���]? �SKD��S �T���{�       ��w hj,a� �pႧ�      `�9r�]? �c� g���w      `���� �T� Ў/       ,�a���  2�̴$ m8�      ���� M�Rk�� m8�      ���� M���w       X2����D�w hÁ       ���֖�~ hǂ; 4�e       �d�����@;Ղ; ��n       X2.\p� ���^       X2��l��y� 0��Z��w       XN�{ ��Kfz� ���        x �d����d��      �rr� ml+�@#ޚ       K�[������
� �@�U�       ��; hf��Z��Os      ���v hf�D��; �1�        <�v ��v	��@+Gz        �j�  0�V� ��z�        �q� �R�J�U� �p�      ��t�w  ��q�Kf*�@
�       �d�y�!"Vz� �)�̭
� І�;       ,���{�z; 4Rk�.q�w �^       X2�i� )�l���� � 3���        �w h�ֺ�� ��Z��f3+�       �D���zg �	�(��; LœO>��       Kdw� Ўw h�S�       �\�qt� ��Z���R�C/       ,w� �Nfn���� �����       K�]? �������t�      �%� ��Pp����;        pp���q-�@K�8>�;       p_��;  LEfn�q7{�����;       p_���R�f����� ��(�      ����f(�@3�8^)�0\� &���       �������X� �b�+e>�+�@;O�;w�D�       ��2ӛ���#G�\)�y�w �����.      ��� moo_)W�\�� ���|�       ��<�;  L���ǯ��l�[�� �T��B�       ���q��� `BƏ>��r��ծQ `Bj���;       ����F� 0!Wg��x��~�k ��_       X�;  Lȕ��Qk��7 L��;       ,��lv$"^� &�v�=3-�@;�{�����!       ��;v셈X� &�v��� ���+W�x�       �0��; L�Ո��K� �}�w        `w��?� &�b���ŎA `r�      `����>��]p��c ��?�        �]f�I� 0%��I�w �"3�]�       ��j�YkUp��j�#n�o~  ڨ������Wz�        ���[o�O�� S���F�(�ߜs �Y�z��7z�        ���� ��8�������|�0       ���o{g ��)�\�Pp�n2S�       �;} h�f��DDd�'}� �$9      ���Zp��J)�F�(���h� �s      �s�ܹ�B� 05[[[��� ��WΞ=�\�       �m׮]���ѭ �Y[[�q�?�W^y�jD\� &hǿ�       �m>���� `�������;�2��S �2w       X �w� �ާ/���Vĝ��t
 �Uku(      �Rk��� `�n��+�@G����lv�w        ����_���z� �	��eWp���?~��z�        "�a�� }�[p��*�@�;        ���� �(J)�       � j�����Z��7�|������u �0�Z��;       L����W2�s �}��n� ���3g��N�       0e�.]�fD� &�V�]� ��Rʷ{�       ����� `��`��Z��w       ���tw �(���qH      �N�y�!"�c� 0U�0|t�Ϸ
�FD� �����_�       ������ӈx�w �����o��V��ԩS�"��.� �\YY�O�C       �e�7�@?�^{�7?��~�a  ]8,      @7�;  Lؿdf��A� ��;       �7��J��۽s �T�Z���
� � j����o?�;       Lɉ'�,"�� �*3���]p�u  ��k׮���!       `J2�ozg �)�����w ��̿�       ��֪� ����� ����       �T�>}����V� 0e{.�g��; ��ܛo��G�C       ��R�KD��� SVkUp�E��g       �Ff�������Qp/�(�@g�       Ќ;z �lς���~���j� �Cf���o���;       <�Μ9�BD�^� 0u�8����(��f�1"��@G��c׮]�v�       �8+���� ����+�\���_��Q `����       g�����  ��]ߩ���~ 4Tk��3       ���ܹs'"�?�� ��]����������9s���       ����������s  (���% ������       �1��� ��Z����� t�0       ��l6+�w�s  �����8~�& ��?�я~���!       �qr�رoEėz�  ""b����ʊw X%3��w       x����� � ���=���܇a�eD�&� �=�R�      ���zg  ~��ѣ�/��:u�Z��7m" ���gϮ�       ���g��^f�a� @DD\����wOo���{DDf��y ���Z����w�s       ��`�� ���̬w�pǂ{��� 8(�k       x2���  ���N?ܱ�ۗ�.�s�����!       `��9s�Z�� ���Tp�%ubǿ�       �܋��C  ���^J�šF ��?�        ���;��������ꢛtUEIL�"(��yf�g��a�e�	K�^�0��#������cB@6�� �YT`�e�Q��FԤ;KwW���c��z��s�����oչ�O���|�I�RzZ� �[x� &���V:       &Q�۽OD<�t �ORJ���8q�#� �j~~~�q�#       `�|�=��  �ɚ�]v�Mq�H� �5�9?�t       L����J7  �b�s���pʁ�I_M �N����m�#       `�,..^�RzH� �[|e�Ν'N����SJ_Y ��n߾��#       `����<#"R� �[�p�/����~ (#����       0a�Y:  �V9�/��k��眿0� `#�����]JG       �$�t:??Z� ��?�N;pO)��C @1ۖ���R:       &AJ��� �Bgڪ�v�^U��; ����       gW�u�RzF� �;�/��k���t�M�� ��z��KG       @������8�t pJk�����#�+#� 6��9���       �f9g! Z(�t�}��z���v��s>�2 (�9�       ����O.� |����SJ�t_?��=�d� ��n����       �F۷obD|W� ��θQ?���l �zv�        h��ҳJ7  ��s��~Ɓ��> ��Rz��C�fKw       @�t:�{F�ϔ�  N-������a ��{�|��O(       mRU�s#q �^���8q⯇� SJ���       �-r�)"�W� 8��`pƍ��_~�?D�ׇZ ��8p��JG       @�z�GF�E�; ��:~뭷�p�o8�����wH1 ��m���٥#       �r��: ��_�u�|�oX���sC� F ����b       6����s��zj� ������Y�9gw h��v�?]:       J:q�Ŀ�9�S� 8���Y��g��� �����W�       J�9?�t pV�}ff�� ��鋋�w)       %t�����(� �Y�y���n����<�" `T�<�^:       JH)�B� ��2p���xD�0�" `dr�/(�        �v�����xN� ��q߾}_;�7�u��s���{ �{`��yD�       ��o����]�; ��Z�&}U����; L���..�        c�� ��[��� 0]�������#       `:��#r�.� ��gW�M�����|fc- ��l=~���KG       �8�K� 0QV�I_��}yy�� &DJ��Çϔ�       �Qj��n�� ��䜇7p��+�_�P 09���~�t       ����m�# �U���/��j�qU��>�� `�RJ�       S���*"~�t �j�ݱc��j�q���Ҫ�� Z�g���}JG       �(���?!"�{q �k٢�z��s��; L��+�       L��`��� ���^U��Z_ P��<xp�t       Ӂ~(���� ��������`�����o���#       `�fffvGD*� �^UU�ޢ�z�w�ޯG���U �s�ź�W���       �f�~��#♥; �59v�ȑ/����:x[��� @+\4??���       0���?E��� ��|�����~��)�O�� ()�|I�       بC��F�ť; �5��Z�yM��� Z�ѽ^�A�#       `#�9�8�t �6kݠ����\[ �9��       �A/.  ��Z7�k��OF�`ME @<���ܳt       �G�4����(� �]UU���۷���� �6�:33��t       �Ӯ� �����ݻ����i��s^ӂ h����u]o+�       k������t �.kޞ�y��R2p��t����疎       ���"b�t �.���y��X� �����-�#       `5���{D�sJw  �s��Z?����̌�; L����J�       X����]��t �>)�5o��<p��K�&"n^�� �v�9_�sN�;       �L�����9�,� �� ����~h���RN)���x �5���W:       ��رcGo&��    IDAT�]Jw  ���}��ݲ��y�1��T< �*�K       ��,--mM)�b� `C>���k��X�� �v��n�a�#       �TN�8�܈�W� `�r��ڜ�k��RZך h�����       ��><�s�S� ؘ�n��5p?z��'#��z> �Ɠ�����       pG7�p�S"�� ��������Għ��Y �5����       �F�9UUui� `þ�w�ޯ����G���x �U���v�S:       ""�����\� ذ�������:�� Ze6"��;       ��s�/� ��X��|���`�w �)��5MsA�       6�^������� �ƥ�ֽ5_����[n���X^���֘��}�#       ���(  �����i#7M�x�F�  Z������.�����t       �O�4���w��  ��{���z?���OZ�� h��[�l�;       ��R�  `h6�1����c�< �9�_X\\�W�       6��i/� �G7���SJ� h�m+++^q      `�RJ��t 0<ݘoh�~�ȑ�Gĉ�� ���^q      `\z�ޣsΏ,� ���L��{]׷Għ6r �*�VVVv��       `s�9�R� `xRJ7^r�%_���GD�?��3 �VyQ�߿w�       �[��y\D<�t 0<�ؖox�zB h�;�KKG       0ݪ���� ������ 8���n�>�#       �N�n��D�CKw  �Պ�/���OG�э� �ʝRJ��t       ӧ��*��˥; ��lݺ��=d��;v���>��s ��������/      �t���{fD<�t 0t�]XX�y��lx�1����֙YYY�KG       0=:4^o��4�M�P�)��� �u����~�t       ��ȑ#Ϗ����  �/���㜡ܫ���a� �N�9�j�       &_]��"�%�; ����a2����]��_�Y @��\�4�*      �d���QD�W� �[�9��a4���I^q�)�Rzi�       &����r��Jw  #󑺮��q�0�CyR h���#;���Jw       0�n��}q�� �h���lXgm��R��� ڧ��n]����8       6����{EĞ� �H�����fgg?ǆu �:���{v�       &�������; ��ɳ��>�Æ6p_XX8��y @+�Z]�甎       `2,..�?"�[� ��ZXX��a6��{DD�yhO� �tﹹ���       L����&"���  F���<l����P� �V����޽t       ���v���Jw  �5��P�+++^p��7_U�KJG       �^9�RjJw  �7�;p���K��R�q�g �s����\T�      �v��z�."R� ��/���O����#"r�2�3�֙����JG       �>u]o��N 6����رce�g}��R�а� Z�i�^��#       h��������t 0zUU���������� 6��s�sN�;       h����e����  �#�����޽{?��� @+=���?�t       �u��:"�R� ��7�|�G�}���)�2�s����u}N�       �j��Gr�;Kw  �R�h]׷�ܡ�#"RJŹ @�䜿~~~W�       ��G�l� `<r�#ٌ�d�>�`s���/����       ���i��/� �O���Gq�H��{��#�Q� �O���-[���t       �W���"�S� ����̇Gq�H�;w�<>����zV�4?]:      �񚛛���  ��S�w���Q<��{DD��C�: h�W�u=��/       h�����qy� `�F�� ���l ��2??���       ������#��� �x��&o�~�-��YD�� @;�;KKK��      �)��t�)� �]����������[SJ�� @k����㗖�       `trΩ��_�n� ����%�\��Q>�.���Gy> �Z��t       �����]D�t� �����Q���G|> �Nۖ����       `����΍�N� ���>�>ҁ�֭[?��� ��RJ?����X�      ��:~��K#��Jw  E����`�����c�g�� h���v��KG       0�~��E�ť; �b�r�޽_�#���1� �P���#���       l\]��`08[J�  e��F���}0��&�R��4���       `c�o����xX� �����z���� ����Q:      �����ߝRzY� ����Ǐhԗ�|�^������ Z�1�nwG�       �'�܉����  �I)���_���g���F�= �n)����Kw       �6�~�'s���t PV����g,����� �ڽgff~�t       �w����`p(���* �^�3p?��>?�� �V��^����       ��7������ @q�WU���h,�;v��?0�� �Vےs�o9�T:      �3����N)�J� ��d��ݷ�㢱�٘���7�� �V��i�c�       �l0���8�t �
��Ec����3�� �vK)u����Kw       pj�^�)�� @;TU5}�ݻw�uD�͸� Z���U�#       �NKKK���t ��p�y�}b\��m��R�r h��6M��      Z����݈�W��oz�;V�u�X���� ���\\\�K�       ���i?_� h�����y�X�'N�x_D�y' �j�ZYYyi�       "�����+"R� �=��z�X��eW\q�7RJ�s�w �wq��yD�      ���رc/I)ݿt �*_صk��y�X�9�?�� @�UUU���N�C       6��i~8���t �:׍�����}' �z�����t      �fT�u�RzUDl-� �K�y���{�D�M� h���K��;      �1���{a���; �ֹ��[n���/��}�Ν'RJ��� @�m����'       �U�4Dį��  Z�u]�:�KKȮ/t/ �b9�Gn߾�E�;       6��sJ)�""�K�  �s��Ľ��E�a������N�sQ�      �i����S��q�; �v�9_W��"�={�|)">S�n ��r��TUuu]ץ~      `�-..^�s>P� h���߿��%..6�9���� @�=|���/*      0�r�i0����- @;圯-uwɁ���� گ��+;��E�;       �M�׻8���� @�]W��b�m۶�QD-u? �n9�s������b?�       L����#��; �V�e�֭*uy�����±���R� ��۷oQ�      �i�sN+++�����- @����ֻ��/�^[�~ �媪����\T�      `����D�cKw  �w]�ˋ�SJ\� h���9UU]]�u�_�      �X���术,� �����K�_t(�gϞ/E�'K6  ��۷oQ�      �I�sN+++�����- @���e�]vcɀ6����� @�UUue�����       ��i�G�cKw  �R��tC�{J�J7  �s>'���C�͖n      �����O)��t 0r�זn(>p?r�ȟE��Jw  �!7�|�KJG       L�C�ͮ���6"�\� �7����tD�{]׃��Kw  �!���^��S�;       ���ѣ�?Q� ��޹s����UU��t 01��_�����!       m��t�s�[� �(ו�h��}vv���8^� �����[:      ��<8WU��1S� ��-[���tDDK�7GćJw  �#��������       ms뭷�����  &��.�䒯���h��=""���� �dI)�rii�{Kw       �E�4OJ)=�t 0q~�t�7�f�e˖k""��  &�=�?���       mp����� X���~�t�7�f�k׮/F��,� L�'v��痎       ()眪�zeD|O� `����ݻ?]:�Z3p��H)�f� L��үw:��Jw       ��4�SJO(� L��������^� �H۫�zm]�[J�       �[��@UUJw  ����V=Rު��ɧ�?W� �H������       �T����`�Ɯ�9�[ ����]�v}�t��j��R��t 0�.�v��)      0.���K��� ��z{J)�������A��� &J�Rz}�ӹg�      �Qk��9�/� L��R�ۭ��ݻ�#�� �ĺGJ�59�T:      `Tz���q�t 0Ѿq�ȑ���v����rJ��; �ɕR��^�wI�      �Q��zK����ݥ[ �������KG|���#"�A랺 &΁n����       �6??�҈xx� `���Z��n����.����z� `�ͦ�ް��tn�      �a��z�<缷t 0�9r佥#N���;v�D�;Kw  �ǏE�      �a�v�w�9�!"fJ�  �꺾�tĩ�r��sn�� ��yz��{N�      ���9���oGĽJ�  �/��ڭvk�[�n�È8R� �|9��l��Kw       �W�����t 0����^W:�tZ;p_XX8�� �(�#�u]o+      �V�^�"�WKw  S�=7��8���#"rέ}� �8?>??�T:      `-����s�o��;�n �CJ���V��9�wE��; ��s��^����       �Q�uUU��DĽK�  Scevv���#Τ�����G#�}�; ��s��N��Jw       ��������Jw  S�CW:�LZ=p���9��	| `�l������ҹ�C       N���=:�tE� `�L�6�����;"b�t 0U.:~��+KG       �J��;?��战)� L����rM鈳i��}�޽_��?.� L�MӼ�t      ��u}���["�n�[ ����.����g����Io)  L�^��yD�      �o���k"⡥; ������1)��q�t 0uf��zS�4^>       ��v�;"�_� FaPU�[KG��D���������Jw  S���x��ÇgJ�       �W�ӹ(���� �����ݻ�\:b5&b�QU�D<� L���x㍗��       6�n������GĹ�[ ��s~s�՚������5q[� `j�M�<�t      ����^?Z� �Z'N�8����51�����#�Jw  Sk&"~���ܷt      �yt��}�� �T{�W\���51���T:  �jw�����nw{�      `��z�G��^V� �z������ѣG����Jw  S�)���S�      `z5MsA�����t 0�RJ����w~g鎵���{]׷G�5�; ����i���       �S�߿sJ��q��- �t�9��_�£�;�b��'M�� �dJ)��i��-�      L��s��9?�t 0�RJ������ѣG�_-� L�*"���t�[:      ��^o_D<�t �)�������#�j��u]/G�[Kw  ��]��z{���^:      �|�n�1�� ��Rz���±�k5q����`0qO� �)���S�      `r-..^�RzSD̔n 6���\O��}߾}_,� lOn�fo�      `2���;��E��J�  ��ߞ��,�9pO)�8\� �<RJ/o��gKw       �%���kr�.� l*oٱc�J���ȁ{D�`0��'���UE������J�       ����$"�^� �\RJo,ݰ^�t�F4M����� ���'N<���/���!      @�5M��xKL�C� �D�aϞ=�I)��!�1�?8�n�  `������߭�zK�      ��z�ޏG��b�7Z ��I)�qR�����`0xCDL�� ��z���\�t      �N�N�9�wD���- ��RzS醍������?�s�X� `Szq�4/(      �K]�۪��&"�/� l>9���{��O��؈��GDTU5ѿa  L�_�v��)      �C�9���]-� lN)�חnب����̼!"�Kw  �Җ������J�       �5M����� ��5H)�N鈍����%�\�՜���  6�s���7Ms��!      @9�^�))�_*� lj�ٳgϗJGl���#"RJ�)�  lj?o���N�C      ���t:���ED*� l^9�K7�T܏=����� ��������,      ����⽪�zG����- ��v����;JG�T��>�Rzs� `s�9?�i���       ƣ��n�J�  �ޛv��}[�a���{D����kJ7  DD����\�      `�><�Rz}����[  ����-����������� ��������n���C      �ѹ��#�I�;  "�3�w��H�a����I�-  �s>'�t���Ⅵ[      ��k�fD��t @DD�����4U���"�D� �������W^y�]K�       �����W��  8iy˖-�/1LS5p߷o��RJז�  ��H)�vv�������[      ���t:��9�.�lw L�w�ڵ������Akڞ� &ޣ�?�ڜs*      �_�߿_J�m��t �7���.�0lS7p?z��"�oKw  ���{��KKG       ��4����u)��-� pߘ��}W�a���{]����  �抦i^P:      X�~��xgDܯt ���ް��p�tǰM��=""����  ������X:      X�Ç��7F�O�n 8��K��T���������Kw  |���xS�����!      ���x㍋��  ���={�|�t�(L��="b0��t ���9�3�i���-      ��u��}���  ��s~u�Q�ځ����#�X� �S�WD����޽t      �z�޳RJJw  �Ɖ�[���tĨL��}����,� p���u�����!      �?�v�?�s~MD��-  ��Rz����ߕ����GD䜯.�  p?q�m�]�����t      ��v�R�݈�R� ��.0JS=p��[������  8�G?~�꺮���2      h�~����ҵ��t �|mnn���4�C����#���;  �����#      `�Z\\�p0\�]� �,^�s���#Fi������Kw  �I�y�i��\�      6��i�r]Dܻt �Y��`����6�����>"�_� `~�i���      �����������-  g�Rz������tǨM�����*  �JW�z����      �iW���fff�)� �9�C��aS܏=zMD|�t �*T9��7M���!      0�꺮���~'"_� `������;KG�æ��u��.� �Jw���v:��     �i477׏��;  ���;w�<Q:b6��="byy���R� `�έ���~���!      0M��������  k�����ۥ#�e��/��#��  kp��`�����K�      �4�v��D�/��  X�?8���6��=""�t�t ���������{�     �I�4�RJ��  k��6Лj�~�ȑ�k�)    IDATk#⋥;  ��~+++�ꪫ�Q:      &Q��{ND�FD��-  k�R����Ͽ�t�8m��{]׃�ҫJw  ��-//_�W޵t      L��i��s���d[) `:��رc�t�8m��VVV~;"N��  X����^{�����!      0	��y|D�1"��n X�+++W���M7p߿��F�5�;  ��n��w�u��t      �Y��{t������-  ��{�^z�WJG�ۦ�GD���n  ؀1??����%�G      �B��}X�����p 0�rΛr�J��sN�^��[  �+��{G��Q��r�      h�N��cUU�?"�Z� `�zϞ=?�RʥC�m������ L��󿙛�{u]כ�g:      �v�~��UU��0n &\J�o�q{�&�GDTU��ҭ�;  6��sss��9oʿ�      ���t.�G���n ؠc����S:��M;pߵk�?����  ��5MӔ�      �R������zDܫt �^XX����lځ{DDUU�J7  CJiw�4��      0n�����D�y�[  �!��[�JJ�Jk�����;  �dq�޽�KG      �8,..^���򁈸�t ����޽{T:��M���I���ٻ�/�����O�ܐLO�FQ�$�"
."����*G����u�kV/Qp����$HB2=���Cý�������g/P���\�u�W�EDP =q����\?]�I�$�������<�ӧN�W�?�  g�A��     ��;��666~;���v9��m��w��uCD�fw  �EG��(;      6�����:��oF�C�[  ΢�;���ڶ�8p�ֈxsv ��TJ��     @5Ms�����.� -Sk}ݝ��mm��#":��JDL�;  β���h�      gK�4Fć¸ h��;v\�1�#���}""ޗ� p��RzF�      ��q; �f���<x�ϳ;�����j��d7  l#w      f�q; �v�[�;��i�4��"�;�;  6C�ui~~���      ��q; ���`0�a���_���  ���;      �fyy����a� �X)e)�a����N���� ��RJ�5M���      �j����icc�7#��� �M�׫����1M���^�w��z<� `�]�4͡�      �+M�|�d2�@D|sv �f���z8ޞ�1Mܿ�d2�>"ֲ;  6�Ѧi~>;      �����y��߈�Gg�  l��Z�k�#�����XXX��R�;�;  6Y��W�F���     ����t����{J)�"� `��СC�1mܿ�Z�Rv ��R�2�$;      �?�s2�����n �
�N�U�����+�����  �;k��h��_g�      �}�Z����k#�G�[  ��o�z�?Ȏ�F�w��rMv �9'"��cǎ}Wv      �����RD<'� `�*�������Έ�%� `��WJ�OM�|[v      ��x<���zqv ���.xOvĴ2p���p="���  �*�����6Msav      �C�4/����  �b��۷o#;bZ�ߍӧO��۲;  ��C#�W_}��g�      �nM�<;"��;  ���n����if�~7�9�Z��  [�[���?p�UW= ;     �v�F�>"�%� `+�R�|����gwL3��b2�,GD��  �b߱s��_�F{�C      h��h�C���GD7� `��Z�u������XXX�xD| �  �J)7?~|gv      �p�ر��t:��-  	�7�4;b����k�  ����'O����iH      ����Gu:���Z��n Hb�|��@��4M�ǥ�Ge�  d(�\���/��      `6-..>����ND\�� ��c�~�q���2�\p?w~�F�  Yj�GF�с�      f����y�n��ø ��J)W���3t�y��PJ�9�  K)ey<?3�     ��q���kkk��n H�竫��̎��gh����k�+�  �:����yRv      ӯ�Zn����G�S�[  �����zvĬ0p�j�������  Ht��x����C      �n��x���3�  ������bv�,1p����o�s� ��=pcc�����     `:���D�|v �����ʎ�%���JD�� ��C��������     �t�����zmv ��mmm�xvĬ1p����������� �)𘍍�w�����     `:4M�k�7FD7� `
��K.���Yc�~�"b=; `
<ymm������J     �m�i�GGĻ#�~�-  S�����Jv�,2D�����""ޑ� 0%~b�޽WfG      �gqq�!�x@v �������7gG�"�{��r4"jv �4��.4M��      �����y�n��#��� �)Q;��8;bV��K�~�c��fw  L���i��     ��������ߙ� 0-J)���z��1����d���  0E:q�x<���      �ƞ={V"���  S�Xv�,3p�����sD�^v �9����G�� ;     ���4��R��� �)�[�~�w�#f���}TJi�  ��7�ر�7�=�5�!      l��i����  �6����Yg�~����j��O�;  �̣���/���!      �]ǎ���xK� |�?��z��1�|ɼ����$"��;  �M)��sss^�     h���Ňt:��DĞ� �iSJ9VJ������,ؽ{�["�/�;  ��K���E�      �w�]w�\��}_D<4� `
�277wcvD����ֺ�� 0�j�׌����      �����o����xlv �4��6���?����g��ݻ_���  �B�Z�ۖ���     ���w��q���ew  L��=��sߘ��gɁn-���  �R{'��{F�у�C      �g��y~���� �)v�E]t2;�-�ϢZk>�  _�7�R~m8��     ��9v��S#��� �)��n����&�g�`0�l����  S�����\k-�!      ܽ���Gu:�#bGv ��*�,<x���mb�~��ZG�����  �b�g�4/ˎ      �]y����xoD�?� `�ݺ���z�Yf�~�:t�"�w ��QJ���h�ew      ��VVVv�ڵ��� �iVk��ȑ#���h�M������;  �X)��aii�{�C      �b�O��6"��� 0�n�v�WgG����&����;  ���&�ɻ�     ��k��ŵ��ew  L�Z뵽^�o�;���}�t�ݫ�w ���������     �yRD4�  3���ݻ�Ɏh+�Mr���OEě�;  f����^�     ��5Msa��]�+� `ڕR�=p��g�;���}�R�F��  3�9��xv     �v���tND����u�-  3ඝ;w.gG����&�����+�  g��z�����gw      l'��2�L���n ���W�޾��7����U��� 0vN&������!      ��x<^�����  ��M&��숶3p�d������  3��k����f�      �ݱcǞWdw  ̊Z�����:���ܷ��ӧ�W� ������^�     �f�����N�ƈ�f�  ̈�w���z�0p�w^q��� ��S��     �F���{k��g�  ̊Z���Tv�v`�Ej������  ���z�i���      h��p��v�o��o�n �!�O&�qv�va�E��M��� �ҍ��.--=";     �-���^�Gv �,)��faa�/�;��-��t^��  3����W���     �Y�4�3"��� �s����(;b;1p�B�^��ַew  ̘~�ԩ7dG      ̲�x�ȈxSD�� ��:�۷����v��W� �}MӼ$;     `�F�=��wE�y�-  3掍��c�ۍ����z����;  fШi�'eG      ̚R����� �YSJy��������n��R.W� ���h���     �Y1�/�����  �A�J)G�#�#��~��"���  3补�_>q�D7;     `�---}O�u�� 0�J)W�z�OfwlG�I:��0"New  ̠'�t�M/ώ      �fKKK�L&7F��� ��RJ��]�'��z�,���  �E��K�����     �i4;o���e�  ̨c�^�o�#�+�D��WF�jv �*�����g�      L������R��� 0�j����ظ6�c;3pO4>[k�:� `F=`cc�]KKK�d�      L��h�Cqiv ��*��baa��D��&�ɨ���� ���Z�5�      ���ѣ�R��� �uӮ]�^����'���� �YUk}�h4���     �L+++�w������ �YUk}�������ܧ�m��vmD��� �YUJ��رcߕ�     �emm����� ��g��v�/eG`�>������� �v�N�s������C      �Z�4?���  �q�����ܧ�޽{��3� `�=bcc��      [iyy�Q�� ���~���������ؿ��xYv ��{�x<�(;     `+���mll�-"�d�  ̸KK)5;��g�>EN�<����Xv �,�������;      6����rD|gv ����`0xv������Z�+�  ���Z덋��{�C      6�x<~fD<?� `�u:�˲�b�Sf~~�=��  3�[���Jv     �f����Z_�� �����>��3p�N��  Z�9M��tv     ��4w�Z9"�� 0�j)��|9�)4~+"~3� ��o��۲#      Ζ�{�^O��  h����fG��ܧT��95� `��Eĉ�px��     ��j<?��:�� �����2�)��������� �x������     ��b4=������ ��J)o���W��[__?��  -p�i�ˎ      �7��a���ֈ��� �8�Ȏ��O�����G��  -P"�������     �{jnn�pD�Pv @K,���[�#�k�S���\�ew  ���"���pGv     ��ZZZ���fw  �A��3���ǲ;�{�S���}�ֺ�� ����gϞ_��      8�����L&7F��� �6(�>�����L&���tv @�R.��O��      �j&��#�a�  -��{��.;����},,,��R^�� ��Z�/---=0;     �4M��Z���  h�Rʡ�������3p����#�gw  ��7M&��     ������#b)� �-j����������ψ}��m�Zgw  ��3���#      ���p�cccㆈ؛� �����#8s�3d~~��#��  mQk}����ò;      ��޽{/��'dw  ���^��#8s�3��2�� �������_:q�D7;     �i���Z/��  h��#���3�3���,"~)� �E�t�M7y�
     H5��D��"bgv @[�R���M��3�3���\ZJ��� ��(���i����      ��N�����  h�Z�gN�>����=g�>�z��''��rv @�쬵�����9�!     ���4��Z��� �&�N���Bv�����:��s�F�_ew  �E)�Q��įv    �-����u�(�-  -�񹹹�fGp��Ϩ�.��dD�<� �e^4�$;     �j�emm����-  mRJ9������;�3�.x]D�qv @��Z�F�у�C     ��[ZZz~D�hv @��Z?���ߛ���g�>���۷QJ9�� �2.�ώ      �mii���c�  -S��� ;����}����_�����  h��F?�     ��p8�1�Ln���� �6�������Av���{L&����dw  �I)����ew      �gϞ�"�_fw  ���˲#���[�СC�o���� ��ٻ����Zk�     ��رc�YJ�$� ���7eGp���D�۽���w�  -�䥥�fG      �0wu:�_����-  mRk������������z���.ew  �M������ó;     ��777�҈��� ��)�\r���/dwpv��H�ӹ2"<�  pv�M&���Cߝ    �{m<?."�;  Z�/���7eGp��H��;G�;  ڦ��}sssew      �i8�bD��n h�:�L^�o߾�����o��~8� �mJ)G�;�-�     �왛�{YD<&� ��n8t��ogGpv��Ӌ"b=; �Mj��v:�7�8q���     ̎�x������  h����#8��[h~~���Z_�� �BO���_�     ̆���ݵַD��� �z����_fGp���T�۽,">�� �6��+���#�;     �鷶�6���� �B�s׮]��l����z[Jfw  �M���Z�O�8��n     �ױcǾ+"��  mTJ����wdw�9�[����MD|,� ���p�-��$;     �N+++�;��["bgv @}����Zv�������۷/���� �6��+��ytv     0}���.��o��  h�����gG���[n0|$"~%� ��vG�N�8��     ��h4�����  h�k>���2p�����K)�� �B�{��7Ȏ      ��p8�UJyCD8� p�}z}}��l>�m����7�Z�;  ڨ�r����ó;     �|{��=ߞ� �F��Ç�Bv���}��t:����� ��������~]v     �kqq�[k���;  Z꣫��oɎ`k�o�^�T)e>� ��J)O�����      r��N��}}D�/� ��j����p8�ak�o#�~����� �6��^=���     l��{�� "��� �Ro����/�l����#  Z�A1Ύ      �����Cj�Wdw  ��j�۽4;��e�����gw  �Q)�Y���G�;     ���cǎ�#���  -��~*;��e�u��a��3�  mTk}�u�]7��     l��h�����;  Z��v�zUv[��}:x���K)�ew  �ԅ�N��<;     �\W]u�J)�dw  �؋8pGv[��}�:y���#�fw  �ԁ�i�;;     �<;w�l"��;  Z��`0xv9ܷ��p8��D�Fv @u#�Ǐߙ     �}���"�g�;  Zj�����#�cྍ���R���  h���z뭃�     ��ZZZ:���(�-  -��^������os���E�?  �������Gew      gO��e�� ���o'O�t�y�3p��Vk��q  �����_]ku�     Z`<?�����  h�I��y�p8\�!��;1??����� �6*�|�4���      ��pة�^;�[  Z�5�^���#�g�NDDt�ݗD���  mTJ5M��     ��777����  -��ӧO_��t0p'""z��'"�� ��zP����     �޹��+���  h���#G>��t0p��<y�hD�iv @�R�7����     �s�v�G��Z 6A����~�m�Lw��p8\�t:Ϗ��� �B�R���p�#;     8sM�<)"~&� ���J)�/�خ���"�^�å��gw  {+�    IDAT��c������     ���y��UQ�[  Z��`0������;_����"���  mTJy����C�;     ��nϞ=#��  -���'O^���1p��\|�ş.�\�� �R�u��&;     �{����R�/dw  �U)�%��������;_����#���;  Z�'���fG      w��zuD�ew  �ԍ�~�}�L'w���p8���� �6���zeeewv     �嚦yZD<#� ��n�t:�����;wi~~���R���  h�o9}�� ;     �bw�Y��  h��z��'�#�^�ܭ����"� �MPk�tyy���     ��v�w\���  h��^p��/s�ܹ[���@  l�s��ׯˎ      �����#J)��  -5)��h߾}�!L7w��~�c��}�  mTJyz�4?��     DL&��#�~�  -��~��{�L?w�H��}ID���  h�奥�s�#     `;k���� ����������w�H���DD\�� �R�L&�;    �$���~�dw  �؋>���f��;g��ɓMD|4� ��7Msav     lGsss�"⛳;  Z���`���f��;gl8��R~."Ng�  ��9��     �����C#�Pv @K�͎;^��l1p������qv @K���h��     ��t��&"�dw  ����/�����w�]�vk��� �F��W���     �;v��"b_v @K��~�Cv����{���wD��E�$� ���}�޽�ˎ     ����N�sMD�� �����>��R�C�=��+������  h�Z�W^y僲;     ����ݻ?"�� �RG<����&w�]�v-D�-�  -��ݻw�#     ������Z/��  h��r�\���2p�^;p������gw  �Q�����;�;     ��v��uyD|mv @�u:��۷o�Fv��������/"ޞ� �B�R���     �6M�<�ֺ?� ��J)W�z�?��`��s6���Ύ  h�'���gfG     @��R�#bgv @�����bv�����l0|�����  h�Z��p8<7�     ڠi���>5� ��&����õ�f��;gE�߿!"ޛ� �B�����#     `�---��� �6��^���'��v0p�Y__qD�fw  �M)eaii雲;     `��Z{�� ����=�ܗeG��5����zIv @��ZϝL&���     �Y5�\k=�� �Bu2��袋Nf���U��v���� ���i�     3��8/; ���t�СdG�.�U��p����܈�=� �e:�dG     ��i���J)?�� �Bu���Av�c��Y�����R��  -����G�#     `��Z��#� �mJ)/:r���;hw6����bD�av @��Z��Ǐ���     �Y0����#�  -��~��������M1�#�yq:� �e�uuu�y�     0��a�ֺ�� �B�ݱc��#h/w6�`0�hD\�� �6���ѣG�&�     �ٞ={����  h�R�/���Ogw�^�l��'O�����  mRJ��;v��     �i���tN)���  -��~��+����;�j8��R��g�  ���M�\�     �h2��G���  -󩵵�gG�~�l��`�?j��gw  ���J)WfG     ���F��Av @��Z/��K�&���3pgK�v�m��� �6����h4zBv     L�R�+#bov @˼i~~�W�#�����p����܈8�� �"��2����     �M�<:"��� �2�<}�t?;�����-�����4� �e��4͏eG     ��X���  -R;��s�9���w��ɓ'������  h�R�����wfw     @��h�C�� ��9����Svۋ�;[j8Nj�ω��� �����՟ˎ     �,��RJ9�� �2���q(;������~��O{��>�&� �E���<�5��Og�     �V;���CD��  h�I��y�����e�����N�^���Z�'+  Ξo��    `�;j��� �6)���z�gw�=����R���s#�s�-  mQJ9t�W>(�     �����s#�۲;  Z�㥔K�#ؾ�I���>Yk�gw  ���w��u(;     �����9qiv @�L"⹽^�Tvۗ�;�����TJ��� �90��ώ     �����qqD<4� �E���dG�������\�� �����fG     �f[^^�)e�� ���?9y��˳;���t�TD�8� �-j��qyy�Q�     ��666�D��;  Zb�����px{v�3���#�W�;  Z����qyv     l���Ň�R^�� ���+����w��#���  -���x���     �����j��fw  �����]������1>���  h�Rk�";     ζ�x�Ȉ���  -q{��y����Og��?0pg��w�Rސ� �?�4�S�#     �l���2"vdw  �A)e����(��)w��d2yID|<� �%�����     8����ED<3� �%�����ώ�/e��ԙ�������LDx� �{���ҏgG     ��0�L���]  �Z�gv����RJ�n�/e��T��z��gw  �A����p�V     fZ�4O����  h�N��܋/������3�N�<yeD|(� ��w�ޟȎ     ����zEv @K����7;;Sk8NJ)?��n �u�֗��    ��j��)�����  h�O�s�9��pwܙj�~��Rʁ� �xĞ={~:;     �R�K�  Z�t�����.��dv�w�^�߿���� �YWJy�p8ܕ�     �D�4?\k�W�  �����^�������3N�>��)� `�]877���     ����  �����^xa��g����p���/Dĳ"b#� `�]����;;     ��x<���=�  3��֟޷o�&3����1>RJ9�� 0�ο�;��     _M���Z/��  h����#�Lu���x����]�v=-"�� 0�J)�{����}�C��[     ஜw�yό���  ���z������pO���L��N�Yq2� `�}������     �+��Sk}iv ���e}}�@v�S�̜^���R� � `��Z�\w�us�     ��ٳg_D<6� `�Mj�?s�ȑ�e��=e��L����#��  ����u�N�zav     |�'Nt#��;  fܕ���ʎ�{���Y����Tv �;����7;     ��[n��'K)���  �aݻw���po�3���g'��s"�f�  ̨�ر�@v     ��'Ntk��ew  ̰�666~j�����C��2pg�:t���k�;  fU�����r^v     DD�|��ϊ�o��  �U�փ������������� 0�������     8q�D7"�dw  ̪Z�;���_�����;3o8�^J��X�n �Q�뮻n.;    ����o��� �+�������gw��`�N+���?+�\�� 0�t�ԩ��     l_���� �[�'��O�z������� g�>��?|�S���"��-  3�O�ӯ{��߿�    ��s�y�=3"^�� 0����OdG���;�r�9�0"�4� `}�d2ynv     �S���v ���������:U]Y*pw� �>�F�#���b �Y��Ą- �@C�:�{���+KHwWUk�3y0����G7��AŇ���"�MY�>tU׹��s#f饪>gy>��ׯ�s��u���^o5;���;e߾}�N��'">�� 0������ʎ     `�����@D|Gv ��hD<��R�C`+�3q���j�K�  c��ʎ     `��� �k��h���C`��3�����J)���  C��m;�    �t8t�Г"�q�  㦔�����dw�v0pgbu:�gG��;  �I��a���7dw     0fff^��  0nj�o���n���b���Z\\�l�ӹ."ֳ[  �I)�Gڶ���     `�>|������  '��O�����ٳ���������v�Qk��� �1��w�S�#     �l���n  3���<{������T�`��Z�����#�� �qQk}�cǾ�m�av     �gee�j�o��  3�5Ms ;��ܙx��:77�����% ��TJy��ݻ���     `2�×d7  ��w�޽�ǲ#`'�3>��t����� �qQk}I۶�     �R����.�\�� 0F>{��ݻ�;�X����v����  #�:??iv     �e8�n  '���4Msgv�w��`0����  㢔�#�     L��~sD\�� 0.J)k�~�u���ܙ*m�gggo���g�  ���\^^���     L����~ث  ��w=ztv�4L��n���qcD�� �1�c    �3v�С���ސ� 0&���{ڶ�Bv�4w�R�4o���dw  ��K:���     ��N�Ӎ���;  �A�u����ߟ�ܙZ��-��  c��Rz�     ���n��A�� �qPk���~��; ��;Sk�޽�����Z?�� 0�J)�9r��     ��]�v�0"�� 0�lff�%tL5w�����?�E�fv �������fG     0~ڶ=����� �1�Z�U�n���!���������RJ��� �QWJy����Wew     0^�;�gG��fw  ��aD����?���!"����K)���  e��s�?���     ��w�1��  c��MӼ!;F��;DD)������� p?J)�<�;�    ���}hOD|cv ��{�����fG��0p�{8p�3����|v �������fG     0J)Mv �������u{�����Qa�_dii��J)�F ���n۶s�     ����Ջj��:� `�m���>�����D�׻="�Kv �������#     m��pv �(��v���~?�F��;܋�`�/"ޙ� 0��m���     �^-//?&"�� 0�~���*;F�A
܋�m?��t�����[  FQ)����fw     0���  ��������0���>t�ݿ*�<#"jv �(*�t�     =�������;  F� "�ZXX�;;F��;܏^����֕� �������fG     0ZJ)7E�lv ��zA�4������c��Zߚ� 0����Bv     �cmm��Z��  �����4��ew��3p�ж�]�v=5">�� 0���v�mˎ     `4?~|oD<(� `��ѣG��0��$�t�M/�\�-  #f�����#     �׶�l���1 �?�陙��ڶ]��q`�'����A��G�;  F�޵���#     �5??�����O �j�/..�Mv�w8M�,�Z�[v ��9}}���     r�R~8� `��i��ʎ�qb����R����� �sS۶��     �X]]�w��� �QRk���`pkv�w8E���?��t�Dı� ��ݻw?%;    ����n  1���xF۶��7�p���j�O���� 0*j���     v����7E�%�  #dPk���[n�Tv�#w8M�~�u��۲;  F�cVVV�    ���ݰA �G����~����W>.�=z����  ��C     ����ꗗR��� 0B^���^�����@۶ù���k���n ��+:��     ��p����  ����=��0���-,,�]J�&"�f�  ��������     �����Y�� ���'N<uϞ=��!0��a4M��֧G�0�  [����n��A�     l�����"�k�;  F��N�s��7�|WvLw�"�~����� ��{vv�Y�     l�}�  #��Rn�v����Ia�[��뵵���� 0^ض��    �	u�С�dw  �������28�-TJ����ƈ�O, `�}������     l�N��� �l�����gw��1p�-�������"��-  �J)7     &���Wew  ${����3۶f���1p�m����WD\��-  ��t�ȑGfG     ��:��"bWv @��gff�r��7ߕ����I�4�mv @�������     �����Y����  H4��^�������Tz��+"�� �,��g���~yv     [�����G��dw  $��~���0��a�R�9��xwv @�Z빵�gew     �e^�  ����^�����t�����7����,"�>�  C��Ew�q�Lv     g�СC�SJytv @�Z�{w����RJ�n�Ig�;`qq�o"����LN ����×fG     pf:�΋�  �|fff�򅅅��C`��i��M����  �Pku�    0�VWW�."���  H0�����_e���0p��4͡���� �O\]]���     N�p8|AD���  �i���MӼ!����;�RJ�t:ώ�?�n �ae8�0;    �S���vVD�Pv @����z��0m�a�u���onn^�n �aO�+_�e�     ���Ǐ__�� ��J)o���id�	�����R�eq,� `��ڵ�Y�     ��d  찿�״m�������z�?��gD�0� `���Z�#     89����-�<:� `�t:����Od���2p�DM��J)���  �A߸�����     N�p8|~v ��R��v����if�ɺ���#��;  vJ)�a    �x�+_�e��=�  ;���z�������R�`0���x{v ������͎     ���ڵ�ٵ�s�;  v�O7Ms$;0p��ж�fgg�RJ�Pv �����ynv     ���Z"�y�  ;����`��;�P������ʣj���e�  l��ݽ{����ݻ�    �?�����xcv ������w.,,|2;�np��������Ԉ��n �f�b0\�    ��+�<?� `�]k�ܸF��;��^������ ��Vku8    0�VVV.��^�� ��6k�����wg� ���;���in����� �͞������     �S���E�lv �6[������s�0�v����Z�[�;  ��=�$     ���o�}WD<;� `��T�4�!;�w�0���ݻ���quD| � `��Z�y�����     ��`0�*"�� ��~w0<?;�o�0�n��OE��qWv �6yPD\�    �?��^ �$�눸�m�����Èk��/:��u��� �J)��     �8r��#K)ߛ� �M��t:�7M���!��3p�1��v�XJY��  �&�:|��Ɏ     �v���Ϗ��� �ND�5�n�=�!�3p�1���Vk��gw  l�R�s�     �����9��� ��PJYh��M���1p�1r�ر����  [�����n��A�     �j8gw  l�Z�r�������3p�1Ҷ�����U��� ��Tk=wvv���    �i�M `B��c��gG ��������ݝN璈�Hv �ۛ     0������Z��;  ���g�m;�N��;��n����pxED�[  �пZ]]}lv�e`    IDAT    ��)�썈�� ��>Xk���m?��:wSKKK�3"�Dĉ� ��2=�    �����Ϊ�>-� `}jss��~��������k����dw  l������ώ     �����D�Wfw  l��Rʵ���vp��a������Z��;  ��y?�    0-j�^� &E-�<����vvpf�a4M�TJ��� ��Pk}~v    �4XYY��R��fw  l�Z�^������3p�	PJ�G�}N)���[  ���:���#     &�p8|nD�� �-������`k�Äh��Ǐ�""�Wv ���t:��    �Fm�ΕR��� p�j�o^
�	b��[n�������� �3����Ύ     �T���WF�Wgw  ��wonn^׶��`��ÄY\\��N�sY)�s�-  g�N��';    `R�R��	 ����R.��������;L�n���Z�3#b�� p��     l�Ç�ˈ��� �3p��rI���pv���aB5M�˵֛�;  ��w���<*;    `�t:��� 0�6"��^����!������.��*� �<;;     `��q�3�֧gw  ����iޔlw�p\p�M���gw  ��Z��������     �w�y�E��� ��Qk}Y�4�)��^�0���ٳy����#��-  ��ˏ?~Ev    ��1;  �4�R�4/Ɏ ���;L��m?733seDܙ� p�     l�����*�\�� p~g0<��R�C��g�Sbqq�o;�Υ��� �SQJ�pee��    �q���������  8E���ظ�m���`g���v�冀^ǲ[  N�LD<#;    `<3;  �}��rɁ>��w�2�~��J)�Eĉ� ��Uk}N��dw     ������Dģ�;  N��"��^����`g����z�ώ��� p���#G�7;    `\�Zo�n  8Y��ϕR.o��}�-��3p�)�4�ϕR~4� �d�C�/     ��m۳�y� `l���{��d� 9�a��z�WD�Ofw  ��k����ώ     7���WEėew  ��ZJy^��}v�����`0�F�k�;  N�������    �qSJ�B& 0j�z��Oew ��aʵm;O��7e�  ��0     �`yy���}�  '������#�|�@�m�>77wMD�iv �xܑ#G�    0.j�7�} 0���`0xQv0|� ���p���ܓ#�/�[  ����泲     �A���R��� � ~{nn�m��C��`��o��G�ǳ[  ��3o���]�     �nyy�����  ��]333W-,,�F��;�O,--} ".��Av �}�������    �1���  �����p������f� ����g����Z��_q �H�.    ��;|��|)��� �������/--�]v0z܁{����7F�0� �^\q뭷~Ev    ���t:�F�y�  _���Z�����v0�܁��4��SJY��  �ssss�fG     ��Z�3�  ��F)��~����`t����뽺ֺ�� p/��     0�n��EĿ��  �5"���vߘ�6w�5M��%� �K<����ߜ    0jv�����	 FO�i��Ɏ F����R��ݻ�o�n �b�N��    �QSk�& 0jV��YɎ ƃ�;pR��ݻ1�)��-� ��R�Ѷ��    �{���|WDx� %?�������0NZ۶���ظ���?�[  �������͎     no F�?TJ��!��0pN��7�|׮]�.���e�  DD�R�     DD۶s�'� �o�����m��!�x1pN����'777/��;�[  "bϫ_���#     ��޽������ ����s�9�)ǳC��c������d8^�� L��>���_�    0�x	 ��wnll\�o߾Av0�܁Ӷ������'G�g�[ ����    �j��z�W�Z/��  ��_��'8p��8m������,�\�m d�����͎     �277w}D�ew  S�#333.--�]v0�܁3���������8�� L�������     Yj���n  �W���q�����d� �����~�ͥ��G�fv 0��     S�ȑ#�,�<:� �Z���>�i��e� ����2�^ﵥ�gGD�n �ҷ���<*;    `��8q�� `:�R>7/_ZZ���`r�[����lD�pv 0�j�q    ��Rk-����  ��F�������e� ����rM����xiv 0�n��;f�#     v���꿉����  ��f)��MӼ!;�<���h��%��� L���y�ߓ    �S�l	 $�����z���L&w`��z�~)����  �K)�a    0ڶ���k�; ��RJY������ &��;�mJ)��.���n �ʞ���s�#     ������#⫳; ����^���L6w`[�ٳgs0<-"ސ� L������     �͋� �{u�4/Ɏ &��;��ڶ]הRޖ� L�:    �D;|��|D\�� L�Z�����`:�;�m�ϭ��_�� L�K�9���    ����t��ew  S�W�;vc۶��`:�;��������0"ޓ� L��O�8quv    �v�^� v�o���]߶��`z�;jaaᓵ�﫵�7� �l��;    �DZ[[��R��gw  �̓��ʅ����!�t1pv\������̅�� `����>4;    `����_�� ��*��~��ʶm���Lw E���h)�	��� `bufgg�ˎ     �^� ���O�8qq��?�L'w M���pD<!"��n &S��!    0Q:���� `b����ƥ���?�L/w U�4w��#�c�- �D��Ç[v    �V�t:7DD��  &ҟmll<��������;�nii�/#��Z�'�[ ��t]v     �zjv  0��?;;{�q;0
܁��4�_D��Għ�[ ��RJ��Z�ی    ��w�Сo��o��  &�_���<ᦛn�xv@��;0B���;����Għ�[ ����+++�Ύ     8S�N��� �V�3".\\\����d������?��^G�[ ����    ��f  �õ�'4Msgv�3pFN����R�E1�n &��m��    [+++�ߐ� L����'���f� |)`$�z�?���#�Xv 0r��~wv    ��R% �U>OZZZ�@v��1pFV�4�O��/d�  ���8�    �R۶�Z�� �D��Z��������b����i���t�ǳ[ ��Vk�Ӷ�lv    ������ވ��� `�}6".������?����v�o���`Dld�  㫔�U�{��ew     ��R�*�3uw��yr�4��@܁����_�Gĉ� `|u:�@    �X��eʫ�; ��UJ�\D\��vߑ�p2܁��4�/�R��� `l]���vVv    �ɺ�eʯ��  �ֱ�pxi�4��p�܁����~6"�G�[ �������'gG     ��N�s]v 0��_k}\������Sa����i~9"�n ��S�     N�=/R>%� ?��7�Z����3��T�c�i������n �K���Ç�gw     <��Ǐ_��  �ί;v�)�~�Xv��0p���������>1"ޟ� �����4;    ��t:�=� �����શm��p�܁�v�M7}|ff梈��� `|�R���     pVWWϩ�^�� ��R��:���m۞�n8���[\\��N����lv 06.Y[[;?;    �lnn^�ew  c�=�N��n�����3e�L�n�����."6�[ ��p������     ����\��  ��Ow:�+]
Lw`b4M�[�fw  㡔rmv    ��Y[[;���� �X،��u�ݿ��*��D��z���;�; ��Wk�xmm���    �/u���'E��/�TJYj��� [���(��z�9�<'"�2� yg���_�    p/��  �¯w��#� [���8���D���� ��Rʵ�     _���o�UJ�,� m��u:�g�Rjv�V3p&R�4\JyEv 0�j����y�    ������ `�m����C ���;0��=��Z�[�; ��v����/Ɏ     �G�֫� ��Vk��~������b�L��m��N���� `t�R��n     ��h�v6".��  FW)�m��W�; ���;0�z�އK){�; ��v������     �{��E�Wfw  #�Z����ٳ���܁����^[k��� `d�}���K�#     :���� �H{Q�4wfG l7w`*�u�Y�"�� �h*�\��     L�;�c&"���  FS)�uM��\v�N0p�����ݵ����� ��K����ώ     �ׇ?���G�Wgw  #��Rʋ�# v��;05���["��; ��t����/Ɏ     ��p8�:� Y�n������b�L����ň�Dv 0zJ)�f7     өm�N)��� `$�n��{Mv�N2p��-����fw  #��Ç�gG     ���������� ��9>33��K)5;`'�S�i�_��_��  F�9�N��    `��ë� ��SJy����{�; v��;0�N�8�dw  ���zUv    0]j�%"���  Fλ�;�C� f� 2���o��IOz�"���- �Hy����#��;�s";    �����]JY��  Fʰ�z����! ��L��`���� `��7??av    0=:���� ����~�o�L-w`j�m;�t:{#b#� ����    ��Pk-�7I �+�|�s�����L��T�v��*��fw  #���o�}Wv    0������  Fʋ���7Ȏ �d�L���>����� `d|�ѣG�    L�R��� �Hys������l���۷oߠ�rsv 0:j��    ��pUv  026"�E� ��� "���/�Rޖ� ��Rʕw�q�Lv    0�����#"�!� �֟l��}� ��� "J)5"~8"6�[ ���5�Ї�;;    �\�/I ��㛛�/ώ � ���zZJ��� `dx    �6�V�A QJ���o�+�`T�|��Ǐ��Oew  #��ZkɎ     &���ʣ"⛳; ���'G�����Qb��En��OE�˲; ����#G�<&;    �<����� `$k��ڶf� �w�/1^���  �y"    �&�d  �J)?����(�`��|��mO�Zo��  ��Z��n     &����R�� ��kff�G�# F��;�����o��_��  �}������    L�R�S� ����7�t�ǳ# F��;�}��6��  �p8�"�    ���˳ �t�۽{���# F��;�}���,��dv ���j�    l��>$"�� �*��߻w�Fv��2p��N綈�Tv ����+++dw     �ovv���(� @�?�v���0�������gK)�fw  �JDx2    8c^� ��aSJ�� ����=z�U��  �C'    �L����O��  R������gG �:w�ж�zD�$� H��#G�<8;    _Ǐ�$"�; �4�333/Ύ � '����bD�Iv �f������    ��*�x) ��kߛ0�NB)��R�� @*�O    �i����wE�E� @�c333/͎ � '����v)����  �\���vVv    0~��'Dă�; �4+����0.�N�p8�G�0� H�{}}���    ���t:^��)Uk�����Jv�81p8�~����_��  r�ZB    ���Z"��  G���񅅅��; Ɖ�;�)*��8"��� �R��F    ��#G�|GD\�� ���G��&;`�����iWgw  )������    `|�C/C��*��ܶ�zv��1p8���Ogw  ;���0
    8�g  )���v9;`���|�ֺ�� �Rʕ�    �x8r��#"�_ew  )^\J�� ������E�'�# ���+++ߔ    ���pxUv ��J)��4͛�; ƕ�;�i������ ө�zYv    0�j�Wd7  )~4; `�������WE�ǲ; ��UJq(    ܯ[o��+"�q� ����^���� ����t����Zgw  ;����?�?�5�    ��:묳.���� `gu:�g7 �;w�3t�ر���  vTgss���    `t�Z�	 ��M�n��� �����m��R�m� ��r8    ܗ���s"��� `g�×e7 Lw�-p����D��; �u��Ç�#    ��Sk�0"�~ S����KKKo�� �� [�m���p�; L�sJ)n`    �/@���������Ia��Ev������� ��rH    �m�v"�� `G�j��}Gv��0p�"{��ݨ��<� �Q��m;�    ����;�q�� ���a3�������🍈�gw  ;�+�9�    ���Z��`���i�?Ύ �$� [hϞ=�����)�
    �b��˳ �SK)/͎ �4� [��ѣ����  vF)��    `4,//KD|Sv �c���z�0i��X۶�Z�[�`z<����ߖ    �����F������;�6h����� `g�R��n����{{����;�]{�$���<I �@[�c�ql��#!m���_Нk�����ԧ��f�S\�pHB�8$�@��!�$���<q�� %�Ȓlyf�Ջ��H������{�^��r�>{-    Z�?e  #��C�});`�A)�F�]� �h�Z�cv    ��رc?o��  F����;�# &��;��\v�eG�; ��+�\s���gw     yz��[� ������Ɏ �T����{��"��� `$J��sv    ��-� �h���۳ &��;�mݺ���; ��px    Sjiii[D�lv 0���?�0���h���gJ)G�; �����i��    �������+� �N���v�!3p�~�o���dw  C�c�Ν7eG     �Wk��# L��8p�� ���`����Nu:�_��  F�!    L�Z뛳 ���ϥ��0��F`yyy)"���  ��?d     �u���+#�� ��}��ɓʎ �� #����݈x{v 0t�9r��    `tz�ޯd7  #q{�4���i`�0"��c���� ��9�   �)��tޒ�  ��O�<��� ���`D������ ��,    ���~���Z���  ���rg�4�ew Lw�ZYYY���d����n{Av    0|333o���� `��YJ����ib�0B�~���[� �Pu�n���    ��u:/:�������}&�`���X�׻="V�; ��r�    �����Z�/fw  C��^�����ic�0b���_��dw  C��i<K    ����>"^�� կ.,,|7;`��$���5� ��o߾���    `xJ)���  �3[�n}[v�42pH077�W��?��  ����%�    �Z�d7  C���������id�����ݝ�  O���    &ԑ#G.��+�; Ŀ+�    IDAT����nw);`Z�$�������|v 04�^\\���    `(�Cv  0<���8p��� ��� ��  ��-�    0�|��	�����n �f� �v���ވx"� �\    0awD�M� �p�Z�r~~����if��h߾}�qOv 0����瞝�    ���R~>"��� G��9�� 0���-//�'�; ���v���͎     �ˍ 0���駟�`v��3pHv뭷~���� �pt:�]    0!j�%"ޜ� ͯ6M��0��Z�����������    �1w�رk"��� �P�XYYqI%@���������  ����Ύ     6����F �P��������� ��d1;  �N��+�    �����Z��z����g������x(� 
�^    0�_�dw  Cq|aa��� �?w�v�;;  �7�u�]?�    lʿ; �T�� ����EN�<������ `�:��7gG     ��t�� ��C��Ev ?`��"M��#�ײ; ��p�    c�i���֟��  ��zwv g3ph��'O�+"��� V)�����ew     �}��=�+� ���:u��# 8��;@�4Ms:"ޞ� ��3g�ܘ    �_����� `(�6M�ώ �l� -����; ��*�8   ���� L��<y�# 8��;@������� `�j����     �����OFĿ��  �MӜΎ �\� -���ߖ�  V)姎;���    `]ޒ  \����� Vg��Rsss�� V�����    `]ޜ  ������>;����X)�׳ ��s    c�i��u:�=� �`���{� 8?w�۲e��Fķ�; ���٥��m�    ���ܹ�Z��� `�=}��'�# 8?w�ۿ��R���  j�����    ��x� &�ۚ��gG p~� -������X��  ���P    ƃoy 0YN����+;�3ph�����#�#� �@9   ��[\\�Ɉ��� ���Zkaa�� \��;�(��-� �+�9ryv    p~�N痳 ���v��5���3p�/"�:� �R�/e7     �Wk�# L��fgg�o ƀ�;�����  `��   @K---m����; ��)�ܓ� ������'O�'"��� F���wH    �̳�>{SD���  �ɝ;w~$;��1pMӜ.��;� �gΜ�>;    8W���# L�Rʯ�۷o9���1p#�^�m���  �!    �P�շ; ��u���Ȏ `��������"�� �`�R�   @�,..�dD�2� ���r�-�̎ `���L)�m� ��\y�ȑ˳#    �p1 L�Z�=� ���;������È��� ``~1;     8��; L�R�#sss��� `}��L)�F�۳; ��qX    -����-"n��  �ײ X?w�1��v�YJ9�� ��6M�5;    �x���]D���  ⩧�~�xv �g�0�8�T���� �@�ڵk���    @Dxq &F)�=MӸ@`���~���� `0j��    �|����� l��;�����8"��� �C3    Hv�ر�Eī�; �������������Z�od7  ��;���    �f�~�E 0!J)��n `������̻J)��; ���v����     Ӭ�j� ��镕��gG �q� c���O�Z?� ؼN���    �4M�5"n��  �w>�tv g�0�:��'� `�Z�{�h    ���ر��E��� `����-��3ps������~9� ش];v����    �R^X�������G�# �w�	��t~3� ؼR�C4    ��� L��g �y� �̙33� ��9D   ����_ZJ��� `�Nmݺ��� l��;�x�[��O�� ����;�,;    �I��-� �@�o���'�# �<w�	QJyGv �y333���     Ӥ��K� ���Z#���0p�����fw  �f�    #r���n���� `��znn�ϲ# w�	QJ�~�
 �ֺ��Z�;    `<��WGďdw  ����  ��`�lٲ�]��� lB)�_;v��    ���=� ��=��t~';��1p� ��r�7#��� ���z���    `��}�� `��Z?0;;��; w�	���=� �oOv     L��ifJ)7dw  �SJ���0� fnn�#�k� �ƕR�4M��5    �ݻw�>"vgw  ��>��`L L�RJ-��3� ؔ�ر���    0�z���� �����R�# ,w�	����ΈX��  6���p    ���rSv �)˵��ʎ `��&��Ç���~2� �8�k    0<M��D�� ��||nn�[� ��;��zwv  �q�֛���?    ��]����; �MyOv  �a,0�N�:��Tv �a�߾}�k�#    `����� �M��֭[?��p�L��i�-��?� ظRʞ�    �D�NgOv �)�ۿ��� ���`��z�wg7  WJq�    ؽ�޻��z}v �q���d7 0<� l~~���Jv �a7?~��    ���ɓo��� ��=z�С�dG 0<� ���;� ��]��c�]�    �ˉ 0��]J�� ��;���ޓL�� `c:���6    �Z�� `�j��e� ��`�:t�"�� `��d    ��h�fkD\�� lا����>;��2p���wg7  v���ǻ�    0	�o�~mD���  6����� ���`
����G��� `C.}�'�Ύ    �I��v�d7  �L���Pv �g�0���N�Z� � ؘ^�wsv    L�Z�� `�>������ ���`z�;;  ذ=�    0��E�u� ������d7 0� S�ԩS_��  ֯�r��޻%�    ����ʛ"�� `C�|��^��� F��`J4M�/��vv �!�N�8���    g��=� ����޽{{� ���;�tyWD�� `C�d    �83p����t\�0E������."�<� ؐ=�    0���y^D�)� ؐ�����uv �c�0eJ)��n  ֯�rý�޻%�    �Ѯ]�����ew  �Wk}Ov �e�0e�{�ߋ�3� ���<q���#    `�Z�d7  ��e˖�eG 0Z� S��[o�ND|4� ؐ=�    0�J)7g7  �?o��ofG 0Z� S��M 0��   ��=z��Z�Ogw  �WJ��� F��`
�޽���O� ���R�o�fkv    ��Z��DĶ� `�N�R>����L�}��-�R>�� �O�u����ߘ�    �ֺ'� ؐ���>����L��e  ���tn�n    �qRJ�M �P�ն`J�L������G�7�; �uۓ     ���ѣ��Z�� ��m۶�Qv 9���޽{{��dw  �SJ��i���    0z�޵�{ ���߿�Lv 9����� `��Z��޽�u�    0J)7d7  ����mZ ���;�;x����� ���Z�   ���� ��ۧO���� ��L�RJ���?� X7�r    pǏ�Fě�; ������i��� ��L�n��I' 3��k�%�    ���_��k#��� `}lY 0p�r���_��  ��w�u׿͎    �6��z	 ��?��%/y(;�\� DD��+ ��n�{cv    ���; ��R��������  ��; ��vߛ�  ���9    ����  ��%� �q���/G��dw  �b�    �q�ر�G�K�; ��+�<>;;��� ����� ��+��ΟȎ    �6���.� �1Sk��RJ��  ��; ���7� X�����    ���`���}�3� |�����"�s� ��8�   �U�� ������Ɏ ����Z�_����ޘ�     ms�ȑ�R^�� �]���� ���; ���t~/"jv �f���;.͎    ���!"Jv �v�nץ� |��; �w�����R�4� X����̛�#    �Mj��g7  ��7���_̎ �=�8K��/b`�ܐ     mRJ�1� X[ �b��Y����#��� ���;    |�ѣG/����; ������ ��������#"���  ��ڦi�fG    @�Z�����(�<2??��� ����s�R>��  ��%�v�z}v    ��`��ZmT 8��; ��v���^v �6�~���    h	w /� �}�8�-���͈��� `mJ)�    �zǏ��Z���  ��K���� ������Y 74M��;    ��c�=vUD\�� �M���� �� �*�| "jv �&�߹s竲#     ��`�t:���n ���X����^k�\v �f�    �j� 0V����|v �d���|(;  X3�w    L�� ����~��R�; h'w Ϋ���� `�n�    �,w�u�+"�'�; �5s�" �e��y���5"�&� X���}��/͎    ��n� 0>�q�ԩ�fG �^� \P���� ����}O0   0�j������`�4�� ������$ ��R��    �ķ1 ����n ������������ew  k�f    �Α#G^���  �䩝;w>�@��pQ��g7  k��cǎ�Hv    �R��ƈ(� ���Z?�o߾�� �����*���x�����Ɏ    �Q*�\��  ��G� h?w .��.{8"��� \\��a    �ƥ 0�۶m�ǳ# h?w .j�޽���� ���);     Feiii[D\�� ��}���?�@���&��g7  krm�43�    0
���WG��; �5�Hv  ����59u��'J)��; ��ڱk׮+�#    `���`<�R�G�# � �I�4�k����  �ġ    S���[ ��G<��� ƃ�; kVk�pv pq�V�z    L�� `<|$; ��a��z|4"z� �E9�   `�;v��#��� ��J).U`��X����oE�g�; ��z�ѣG��    ô��� ���ggg�*���a��z�E- �_���Ύ    �a�t:�f7  Wk�h)�fw 0>�X��e  ����^   �D��^��  ��G� /� �ˡC��_��  .��b�   ��j�f&"���  .��ɓ'?��x1p`�J)��  \ԵM���   ���}���FĎ� �>�4ͳ� �c ֭��?� ����K/����    0�n��� `MlL X7w �mff澈8�� \X��w�   �D��^��  \����ǳ ?� ������Dğdw  �   �	�r h�/,,,<���1p`�<! ��   ��s�m�� "^�� \X��c� �'w 6���},"jv pAW.--�Ύ    �Aڶm�uQ�; ��ry" b���>|�Ɉ�Bv pA����7fG    � �Z��n  .��^~����x2p`3<% ����     �� ����Ͻ{���; O� lX)�SR �r�Vw    &F�4���j! ��M	 f���=������  ί�zm��dw    � �޽�ʈ؝� \Poyy���# _� lX�4���	 �X)�_;v��    0�^ϋ� �~�ַ����# _� l�'� ���:�   `"�R|����%`S�ؔ~������ ���   0A|���+���)� l����7"�� �9�   `�;v�G"�U� �=���O�yv ����M��[ h��wdG    �f�z�k�� ��MӬdG 0���� �@�͔R�Ɏ    ��(�x� �φ�M3p`�v���PD���  .��    c��zmv pa+++�� ��3p`���۷�gw  ��   ��Uk-� �ݗώ `��0(���v�.;     6���~eD<?� � � �������av pA?~�ȑ˳#    `#J)o�n  .����0p` ����>"��� ��C@    �U���� ����t:dG 0��R�_�@��   0�������}&;��`����Z?��  �_����    `���y^D�:� ��Of 09��n�{D��; �ՕR^�4�Lv    �ǎ;���-� ����1p``8�TD|.� X]�u��;���    ��(��!� ���.��G�# �� �'� ��ޘ     �tMv  p~��������� `r�0P�VON@�9   `ܸ� ��V��2p`��m��pD<�� ��s�    ��{�ggD�2� 8����Of7 0Y����������; ��jiii[v    ��3�<����fw  ����Ç���d1p`�j�����ں����    X/@��qv  ������v�� �b�~ߡ     c���[ ��� g����8q⑈�vv p^�d    ��@��z��� �<� \�4�Z맳; ��zcv     \�w�qiD��� `u��/>|��� &��; C��t<A �u�ѣG/Ɏ    �ٲe�"�dw  �uv  �����p�; ��L��{]v    \H��Cv p~�N�6��0p`(<���fv ��R��A    Z�7, h����� �L� E)�F�� ��j�   h;߰ ���r���'�# �L� M)�ST �Rn�   �͎9�xYv ��Z��� L.w ���rv p^����;weG    �j:�� ��\z�0�04�RD|+� XU���^�    ����� �b�N�� &��; CSJ�� h�7f    �jJ)� �^������� &��; CUk�$ ��5�    ��Z��; ���� L6w ����  �   �:w�u׏Eċ�; �ՕR\v�P�0T��bD|+� Xտ>z���#    �_*��1� 8����� �l� U)��Z��  VUz���#    ��\�  ���/,,<��d3p`��  ��a!    m�w h��� �|� ���� ��J)o�n    �����A h�R��; Cg���:t���� `Un�   �5���"�ǲ; �խ��ܟ� ��3p`�J)5"��  Vu���⋲#     "bffƋ� �^_=|��� L>w F�U �^��k�     "��b� �e��H�0�V�� @K94   �-j��U@K�~ 0*� �ġC��6"���  ���   �6����x}v ��Zk�?;��`��(}:;  X�Og    �����#�� ���<??��� ���; #�* h����;";   ����v�4 �e����02�n�?; �R333   HUk}}v p^�g 0=�����GK)�gw  ��:;    ��� �Sw F������~:� 8W��u�    L��� �U���C�����0p`�j��e7  �2p    �ѣG_/��  Ve��H�0R�^�S� ��.����4;   �����\�  -�2C F����ZXXx<"��  �Qfff<   @�R��� ���+++dG 0]����� �B   H�� h��u뭷~';��b�@w h�)�Z    IDAT'��    dq� �P�����3p`�z�ާ� �U�.;    �鳴��;"^�� �����0r� ���Ç���G�; �s\�4��#    �.�>��UQ�; �s�lٲ�� ���; )J)~� �e���WdG    0]:�����>���� Lw R�Z����ݮ�D    F�7) h'� R������5� 8�U�    L��� �s��}w R������_��  ��0   �����{�D�� �9�K)gG 0��HSk�K_ h�Z�U�֒�   �t8y���-� 8�g���NeG 0��H��t��}v/..�<;   ��qUv  ���� �^� ��v�DD��  ���v_��    �Ը:;  8W��0���e�@�[n���hv p�~���,    F��� h�^���lv ����l~� -SJqk    CWk-� h�R������2p U)��� �n�   `�9���� �l�V�����le  �xɑ#G^�   ��s� ���
�f�@���]D�cv p�Z��E    ���� ���ʊ�; ��HWk��� �l�N��"    �� �ϣ�~2;��f�@:O[@���   �as�; ��C� `�@�N��`v p��    �m����Z�e� �9\R@:w ҝ8q���tv p�W5M�=;   �ɴm�6, @�z=�����tMӬD�g�; ��tw��yev    ���j� �������ˎ  w Z���+ h���    �L� �>��K)5� �h�N��+ h���    �L�w h���  ������������ �,   ����m��� �l�w Z���V���;���  �rU�4�o   `�VVV^[�; �(��>q�� �`� @��%0 �ˎK.���dG    0Yz���� ��j��i��� �0p�]��efff^��    �d)�\��  ��f��0p�5j�ED��  ��   ��*��6� 8��; �a�@k���}+"��� �@����    L�Z�� �Yz�^�3� ���h��v1p   ``�=��x~v p��>|��� �g� �J��� ��eKKK��#    ��~߅
 �2��� �_2p�U��u�����    L�R�k� ���Z�n ����V����jD�cv ��V�j   0�5@�t�]w Z���֩��iv p��    �oM �._=p���hw ���  �,   ش�i:�����  ���v Z����)���	 ��5�    ���۷��ֺ=� ��Z�f7 �3p�uv�����x&� ��-..�(;   ����t\�  ����  �a� �ξ}��K)�dw  gyuv     c�7& h��/���/fG �3p��j���n  ���   ���	 ��/����ˎ �f�@+�R<� -��t>��c�~���{����'��!�"*�\�Z�o�1������z�C�F>�-���^�K�J1�����샤1Ɯ�}H�������
�O���]   �=���c�i1>�$)�0UQ 0!   ������Lv ��0U
� Lҋ/���R�f�  n��Zkd�    `5moo?[J��� ��l6Sp`���2) �����O��dv    V�7�  ���Ǐ� �D��)Sp�	���    |^�  ������ �w ��a
 &���   ���� L�0F�,w &�ҥK?,�̳s  7y�   ��r� 2�͌0Y
� LV���K)�g�  n�	   ��}���=ZJy2; p�Ս��ײC �N���Z�/�`:���~#;    �ecc����� ���^x�jv ؉�; ���� �遭��g�C    �Zj�� bl��Sp`���C L�|>�Fv    V��; L��A &M��I�ַ��f)�w�9 ��"���    X9
� 0!��:w &-"j)�g�  ���    �I�U� ��ӧO�2; ܍�; �~� �1   ��������x4; p���  �Qp`��`R�>s�̑�    ���0�  Ӣ���)�0y�/��!; PJ)���g�C    �2�`Z�%;  �F���;q�ąRʛ�9 ��"��    X]�)��t�k�?� �Qp`U�� &b��gg    `5�Z�`:^?y���! `7
� ���  \g�   �e�Z���?�s  ��Z���X	�08d�tX�   `W/���S����9 ��"¸  +A���p�ر�K)��s  ��R�8{��#�!    ���|��� �Qp`%(���{�E��G�9 ��a�ki    �*"��� ��/��Fv X��; +#"~�� ����     L��; LǏ"�f� �e(��J,��t(�   �wH 0FX%
� ��a� `:<N   ���f  n2*��Pp`e�<y�祔�9 �R��K   p��������pv �:�� �w VFD�Rʿe�  J)�;{���    L�0�  ���K/�t>; ,K��U�b ��n�X<�   �i���  LDD��ƨ  �w VJ��G� ���p   �wG 0� �w V��; LG�uV�    ؉�; L�� +E���r��ɷK)��� �Rk�jv    &�8 LD���� `/�X)QK)�7; PJ�H	   ���?x���Dv ��Rʇ/���;�! `/�XE�,�i�j��Ε    ���W�>[J�� ��v V�" ��G� �RJ)������   ����� 0����Qp`��f3�/ ��Z��    �wF 0FX9
� ��'N����6; `�   �;Rp��X,FX9
� ������ @)�֯fg    `Zj�F `>8u�Ի�! `��XU~� +   ������x:; PJ)�z; +I��U�� ��w�    �t�С�K)��9 �R�n +J���4��}e ��o��_�   �4�f3����w V��; +���ӿ,��&; P��Ɔw    ���" �� �*w V�/�`"£%    ��] L���N��uv �<�XY�V_�4x�   �}-;  PJ)��d ��K��Uf� &��;    ��jv  ���Щ `e)����ap�iPp   �|���}����� (e�fg ��K���u�ԩwK)�e�  �S}��   @�����eg  ������� �y)����  �졇z&;    ��� ��?O�8a0�����J��*���Z=^   �� �A������J��gg  J)/   �Wk�Zv ��R�k� �^(��҆ap(�iPp   � L�. +M���v��ɷK)�s  /   Z��+�<TJy<; PJ�u?��  �B������zv �<���3&   @��������� �O>��㷳C ��P> `�E�/� Y����>���    䨵�� L�k}��! �^(���j��eg  J)�x�   h�0�#; PJ)��e �{���:Pp�	��>��   ��n &����� p��Xy�.]z��2�� ������    @w ���Pp`�)������RJy3; �΂;   @Ӟ�  �ťK�~� ; k�� �ς;   @�^~���J)e�  �O���� ; k���Zv �<�ꫯ�   ����?��D�� kA���0�w �w��ŋOf�    `\�� �`�u���Z�w ����<f   4fwB 0�X
� ���'O����~v h]���   � `677-���X�V_"@2��   h�;! ����?�Av ��X�� �<f   4���tv ��L �6�X�V���|~G   А�_~��R�Vv h�Q@ ։�; kcccC� �=���Fv    �q��5��iЙ `m(��6�x�7#�rv h܁���'�C    0��l�~ 0��܂; kC�����s�-j���� Z�X,<j   4b� ����>��g�! �~Qp`��" �E�GM   �FD�� ��z��Cv �_�X7�e  ��;   @#� �$`�(��V�aPp�d�V�]    ���>�� 0�zQp`�9r�R��n@.�]    x��+�le� ��E�w ֊�; k����R���9 �qO�}��   ��u��5C �o8x��g� ��I����gg ��mnmm=�   ��5�͞��  �_����������� �l{{�z   ���� $�	 ֎�; k�뺟dg ��u]�q   `�E�;  HVkՑ `�(��v|� ��q   `�E�3� �u
� �#w �Α#G�,�\�� ��	   ��j�Ogg  �@ ֎�; k����.���� g�   `��9s�K���� и�<�Fv ���XW�P�\u�ܹYv    �G���  ߛ/����� p�)���~�  ���;�<�   ��1��� ��? ֒�; ��! �E�_gg    `��� ��`-)����ap��|V�    ֔q �� �%w ���˗�*�|�� �   `ME�q H6���������Z��~(��4; 4N�   `M�Z���  ����SO�<; �w �V�կ�  �/   �5��+�<ZJ��� ���s�=�� �A��u�W\ �멾�;   ��իW�*; P^�  �E� ���u�w ���C=���!    ����;�� Z�� �3w �����w H6�Ϗeg    ����>�� Zg��u����:u�ԯJ)�s @�f���N   ���� �u]g������ڊ�ZJ��� вZ��    �_q,; 4������� �E����X�D;   �O�Ղ; ���� ���Xk�֟dg ��Yp   X/}�w��'�s @�����Xk� �5/   �5r�С�K)d� ���`�)���f���; ��ʹs�f�!    �?f�ٱ� к�Pp`�)��֎?�A����9 �a�~��'�C    p��c $3���Sp`��r rmnnz�   X�z  �G'N�x/; �'w �^D�r �p,;    �ͱ�  вZ��� `�)���j�� Q�ժ   ��8�  ��� �~Sp`��Z�� Zǲ3    p�3 �\: �=w ֞�; 䪵��    ����~����9 �e: �@�����o}��R��s @�����   ��9�R�Fv h�0
� �=w Z�Fv  hU���W_}�@v    �! ���S�~� ���; ��3 �]�|�+�!    �g
� �("ވ��� ���; ��� ������    ܛ�8�� g��&(��
�< �e�   `����\� 4A��V8�@"�^    �� ��} �	
� 4��ѣo�R��s @�j�ǲ3    poj�� QD(��w �����o�R��� ����'   �
���`)���9 �a����� 0w Z�Kf Hb�   `�:t�/�� d�E��W�C �>h��; �y���    +h6���  ��y �
� 4#"���  ��G�>�   ����  �8w ���@K�  �b�8��   ��'"�eg ���< �w ��u�� $��fV�    VT��� ��y �
� 4�ĉJ)�g� ���ev     >7w ȥ�@3�h� $��   ���� @�߽��Kf� ��(��w �s,;     {w�̙#��?�� ���  0&w �Rk}#; 4��   �jr� �"B���(�Д��U3 ���ٳge�    `o��{2; 4���h��; M��f�j�<1���";    {���  вa���w �r���_F��� Ъ��
   �b�ap� �j��h��; M��~����� Z�u�w   ��t  ��cǎ�� cRp�E�l�<־    V�; ���s�=�� cRp�9��7�3 @�j�־    V�; ȣ� @s�h�w ��1   `�D�; Hb��)�М�l��� �0��   X!�����Xk=�� Z�u�� �Qp�9׮]�Yv h��/   ����a�  �Z�h��; �9}���Rʇ�9 �Q_����   ���w H4��; �Qp�U� ���ѣV�   V��; ��t����C ���h�ϲ @��aPp   X�. ��,"jv ��; M����3 @��~   ��a�� @��I
� 4i� ���   �JQp�$��@��h�l6s�$�Vw   �a�  R�6 �$w �t��U� ���   �
��F)�� ЪZ��; MRp�I����R�G�9 �QV�    V�?��?>ZJ9�� Z5�͌��$w Z�Kg �a�   `D�{ �������� �h�/� �#gΜ9�   �])�@��GD� �hV�Ղ; $���    �]��/�3 @�t h��; ͊���3 @ì   L\D���$�� 4K��f9@�_    ��p  ��> ���@��� RY�   �>w8 ���:�} 4K��f���K�R~�� Zd�   `�j�
� ��h �Rp�i�V���~o   0m}�w��ǳs @�"��'~�� �(�д��K/ �a�   `¶��+�lf� ��Zߊ��� �(�дZ�_z@�    �X,�� @c} 4M���E�[� �Q���?x0;    ;�> �c���)�д���3 $�t���    ؑ�; $�7z Z��@ӆap(�$~s   0Q�Vw7 ���:] ���@�N�<��R��� �(+`    �n  ��; MSp C Ha   `�"�� ���'��gv Ȥ� ��";  �H�   `�j��gg �F���~� ��h^��|v hQ�u_��    ���� @ Pp��u��� ТZ�gg    �O}����B)�Pv h����<w p8�a   `� @��8�� �)��<�����/�Z#;    l>�+�@��0�@��h^�u�(��� Р��|�;�d�    �O�� $Qp w (�w�Y)�7�9 �E�X
   01a� �\�rE���)��u� @����R   ��qg 9>�����e� �l
� p�/� A�u�   �ǝ �8�  �@� �;�  �   `z,�@�| P���RJD���  -��*�   LL�U� r(�@Qp�RJ)���! D��R   ��qg 9j��3 �(�@)e6����  -��   0-}�,�|!; 4�8 w (��r���wJ)Cv h��]   L��֖A ȣ� E� J)����WK)�e� ��D�S   �	���	  �b�x'; L��; ��3 @�>{���    \
� ��ӧO_� S�� 7��W_ � "��    �M�� 9t �w ���; ����)   �tXp�
� p��; �Pk=�� Z4�GS   ���w5 �@g �@� ���� ���:�    QkuW 	"Bg nPp�666�gg �y4   �� �F� nPp�>��R�"; 4H�   `"j�
� �`6����  S�� 7<���ۥ�w�s @�<�   L@��])��� Рz���w�C �T(��-j��3 @�,�   L��Ç�TJ��� ��������  WIDAT�! `*���� � �    0����  �:�  �D� nQk��/ �c7~   @�Z��� �Q�
 p �ED��� t��|$;   @�"�  �� �B� �د� @����x
   �� ��U �[(��sh��0|9;    � ��U �[(��-��C# $��k   �|�0����
 pw �ũS�>)�|�� ZSk�   �� ��A� n�� �� Ƨ�   ��K� �Aۗ/_�Mv �w �M�U� F�eg    ��������� �D� n�u��; ��ϲ    ��W^y��r4; 4HG n�� ������ ZSk}4;   @��� ȡ� �Qp���Z`|P   ��s �CG n�� �� ��    Q�u�g  AD��< �F� n3��; ����3g�d�    h�?�@ ���; ���>sx�V�    ��Z�� @ ���; ܦ��˥���s @kj�V�    ���Vw ���; �ٻ� �AQ   �D�w ߕ_|�w�! `j���|! #��#*   @�Z�� ߯"�f� ��Qp�;Sp��Yp   ��n Ƨ�  w�� w�fg �yD   H�`|
� p
� pg� 0>w   �$�Vw �n ܁�; ܙC$ ��J   @��ﻈx$; 4H7 �@� � ""`|�   lnn>\J�e� ��DĻ� `���>���wK)5; �dw   ������ 	����)���}���av hIDxH   �ax  (���)����s��q=r��9��   ��; ���'N\� S�� ;����� ���|8;   @���  ���  0U
� �3w �l6{4;   @�,���t `
� �� 0���m��    #�� 0>� ؁�; ��:�I YD(�   �lw2 0���I �(��,�����   �ϝ �O' v�� ;p����    F�� )t `
� ���b�0	 �Sp   �; ��= ؙ�; ��ʕ+�Rjv h��T   �����f3w ؁�; ���k����s @Kj�~�   0�3g����� ��z�꯳3 �T)��ݽ�  c-   `D `|WO�>}!; L��; ܝ_���"B�   `D�V�1 0��"�f� ��Rp��Sp�qY   �0�c `|� p
� pw� 0�#gϞ=�   �!�`d�~v �2w ��Z��; ��o�   �Sk�bv hM���� `���.��Sp��E��3    4�] �,"t �.��.,����ax8;   @+��s ��E ��Pp����� Ff�   `<�0�������Sp������� �Q   `$a� Ffl �N� ��ԩS��R.e� ��X   �����677��.�`wV�`DU   �Sk�� �_�p��! `��`��i Q�u+;   @C� ��>��~� S�� ���*���"�j   �x�� ��t `w
� �;�K QDX   ����z��r$; ��_�`w
� �_O��j�
�    #�z��{ YD��� �N� v�u�� �1V   F����pv hM�U v�� ���� �1
�    #�A� FVk�A �](��.f���% �K�   `� F: �w ��b�p��qm�}�
   ��j��`d�`w
 ��Ç;\�����   �Sp��u]��  �Pp�]|�߼TJ�,; ���
   �φa�Bv h�|>Wp�](��r>�  -�����
   ��"� ���>�? �](��"�� 0"��    �/"�E �u���k�! `��`	�Vw ��;   �������q� ��`	
� 0.w   �QXp�q� ��`	�	 #�A�   `�)���t `	
� �� 0:w   ��� Fd\ ��� Kp��qE��U   ��g� Fd\ ��� Kp���)�   �Zk�R��s @K���r�`	]�9d��,�   ���>ZJ�e� �����(����C& �hw   �}t�ڵ��3 @k���r�`	p��Yp   �_�0(��Ȇa�= �%(���?~����� ��   �� ����; ,A� ����av h�1   ���� Fv��� X��; ,ϗ� 0���Ν�e�    XW]�meg ��|����� �
�`y
� 0�x뭷�   ��j�
� 0.� X��; ,�a F����`v   �u�^ `\: �$w X��& ���:��    ����� FTk�9 �%)���"�a F�X,<�   �� 0�� ��Pp��}�  Z�   `�Xp�qu]�s  KRp�%���� Вa<�   �Z��� ВZ�� ,I� ��u݅� ��    ��� �N� ��� K�� ��l   ���� �� X��; ,�a ��   `��Z�fg �����)����a��� Z��   ��ܽ ��j�: �$w X���}M �:�    `�)������9 �%)���^xᅫ��ϲs @C�   ������f���; ,I� �Ɓ FRk��
   �Ν;7���� -�x� ,I� ��Bv  h��;   �>x��,�Dv hȕ��d� �U�� {����Xp   �����] `\� �
� ��V�N IDxh   �����] `\� �
� �7� 0�    �`6��w��[< 썂; �ͅ�  ��    ���z4; ����`o�`o:`<
�    ���:�. 0�Z�1= �w ��N ��V   �}0�{ QD��=Pp�=p��Q��޹   �>�w �� 쁢  ��0� 0�x��Gg�    XCG� @Kj�� �
� ��`\���G�3    �� 0.] �w ؃Z�� Вk׮yl   ���
 ���`o�`��s���f3w   ����z4; �d�X� �(��<xС F�X,�   �Z�; �w �w ؃��ۿ������ Z�u��V   ��,"ܹ ������� V��; �AD�R�'�9 �[   ����  В�����j�r�X� wT�=�����>�%�1,�"q	��
�IHȆ�{2����/R5�}'�]+3��� ���= ��e   �)ܹ @��߿�  A� I�wO (b�;   �� �����p�= �� �� P���   `<w. PGc  Iw ���� �("���    ^��� ��h  I� I��� P$"^͞   ���  Dc  Iw H�;|@�;   �x�\ ��� �$p�$�; ���&   0�� ��J< �	� Ͽ����V   ��>~��� �2�5� $9�@ޏ� ����   0�ϟ?ݷ @!� O� I˲8|@�   �\.w ��1 �$�; ��| �{p   �z��o�Z H�@R�ݿ��HD��   0���� j��=  �� �� P'"<�   ���� �e�; $	� iY�; i���   0PkM� �,��<�; $E�W@���   t>�� P�= ��@Rk�� �xp   �z�Z(  �,��$�; $]�W�; ��   `,��V�]c  Iw H���u��"�w�    ��ܷ @!_��<�; $����| Ա�   `�eY� PKc  Iw Hz���O���� ����
   0�/�@���� I� �8�@���{�   ���< (����/ �$�; l?f�  �߿��
   0��� �Hg�  {#p�z�̞ ��r��   ƹ�  �����:{ ��; l#p�"��Y�   0�� ��k�  �Gw ؠ��
 E�e��
   0H��w �cy l p��eq�"���]   �w- P��< �@� �� u"�w   �q� P��< �@� ��B���|��
   0�� P��< �F� D�C( �^�6�   �Zs� E�E� [��mlp�"6�   �c�; �i�� vI� �����b    ���HD�g�  {$p�m~�  �����   `����� `�� ��� P�w   �A, �R�8 `�; l6�@��p�   0�M� P�� `�; l�{�� ���γg    xAܵ @��� �	�`�; �qv   g�=  ȫ>��= �H  �i� ���[�    �q� ��9{  ��; l��3 �Q�   �r� ��u�@�� 6轿�= Ekͣ+   �8�� �Hz�w H��!p�"6�   � 
	� O� ۼ�=  ��   `(w- P("�1{ ��; l�Z�@�֚GW   �q�� ���� Iw � "�:{ 8�eY<�   �� �Z6�@��+ l#p�:ή    �X&  ���  �F$  ���Hk�<{   �D� �� �$p�m��  �""�    �k�Z��  �F� ��� E�    C�k�Z��>}���! `O� �������tz={ 8�޻GW   �qܵ @���Ƿ�g �=�@җ/_�~�
 ez�~w   �� �XD�6{ ��  $-���3 ��D��W   ��~��Ξ Jg  	w H��Ϟ �D�   0Ʒo�ܳ �: H�@��' �{x   ����= ̡3 ��; $�� �<�   �Z[g�  �3 ��; �9x@���   pss� &�H r� ���	 �z�^   X��= ̡3 ��; �9x@-�    ����3 �A�  A� I���� �Hlp   ����= �q7{  ��; $-�b�	 ��    ��g�, 0�� ��@R�]� �\�   �� ��Z ��@��_ (��   `�eYܳ ��d 9w H��0 ��   `�; ̱,�� � ��Zs� ���   `{, ��k� ���
 y~?��K_   �1�����~8�N���������#�!�� ��˵��?��n    IEND�B`�PK
     Y�#\$�3  3  /   images/7ade412b-fa94-47ea-987a-d6c9baa14438.png�PNG

   IHDR   d   �   {��n   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  �IDATx��]�Uy�f���o�'YB�D��[��Z,� B���c�6E%�S�֧�$��XJ��Q�Z�h}
�<-�#�XD�b�f�Mv�ww��ߙ���3sw���͝9s�ݻ��/{�ܙ3��|�9�s���"��{�,W�\�r�J���[�%�2����,���"Kv���=�����F��t�X�gYǲ�����%΢��X��fy��,a�S�w!�ES�c����.I��Pﰏ��{Y�ay��Y^f�W�W@���K,og���d���_����%I��$���4�����7^����;�2K4x����7n
�1e���d|��f
z�-7��X^a��X�c����D�����3Kd؉DXַ�Ί֌���;X�IV�Hj��,��Ĝ��E:�p,�SD�Q�?G�ߨ}��BѠ�L�rEc-���s��ɸ�,+c�Ҥ����Z,
�5�_��cq�-��i\M�3l��>��Y�H��W��繐���!����(+���NQOG��QT�Ε/�\8����l�Q*&'bl���#�C��̘��g��#�� CC>A2,���d��1����"��%���Y� y�% �шF���ζ�l<�4U���<��_�9�岘�%�#`�*cj�f�}�U��S B\ځ�6�oPiq��^��J	u��{��ՃS~4��@��n�.&�0eu#k0M%��|�D9!K�(�q��5*�"3?ux@Kt�c-�%��~��2ۙ����d͈�d���E�5+���<2��)�9@>�f�X2���Y��D_���:���s4&�
�~2K������ P%��T�e��JG!�� ��5�N]�C�'���͋�'�C����E8/ЄW�)�+��!{5�Q���l�K�͖Q�[�&(Td9������;���yd8@c���k�:�J��>49+���t$��,��H��.��k�� v,H�T�ĩ����F�S�!�y��`�����&e'S�����}�(�د;!'xh5y�X�Z�E��PL'�b��?�B����W`u?VC1p�ɣ�Q�[a �e#/Q��CsB��/�۩ق�`��P����O����k�Q�΁DX���g�E1d\3�E�a�;��+�iё�zӰ!`��F+� Yy��$�p�����鲿x���Me� �`B�|����|�~�򘘩�u%E�9�C\h�k�i*:�p����h<B �eӵ��1Jƣ�4em�O��)�ȭ�lhb� �I��6ߛ��u�Đ��!d��@�������4;����!�Ў<��hV�&���E�o�v�źh�"�/��ά�Z���iJ���E�/�\伣Nh�0W�Y��U�"�@�Y��\�E�/Xl��g��!~`/�����i0��(G�f��1�ri��b�R�o��XX]O��-RO��"���DZ&�a &���ݢE�_訲�İA�4�%ur���ei�%��zb�@���U���r��t�LH�<q��]�dZb/�4[EZ@MD��]1L��J]�R�h��K���N�����7!֬FZ���*Z�@�h��Y�8��_��}b���>>�כ�t6[�Y�l�B��;z�EP��-[�;_@����}������hk>� ���I>�W��-ш�#H�Jщ�b6��du�%��Yv�-Wp�#�9/tXb��q_REK�zXC�wdŦ;hb�gjN5��l`IA3��(���!�͞�V���)t��銑�`��a�!��u�=y�H��J㿤�u!G�w��,�C7�y,#���~A	A�8�a)�Q]h�k�GE��|��tir�B�����.��{,y>�����&\u���$9�y�@l��4]�i�����]�!.s�M���G�wٰ�PGk$��(�Q"���vZ�R��zL���?���gĊu�GGZ��&&R0�J����R9/�Ē2M-�wş�|��kJ.��\O��x�J�#��D�S���l�@��I�ɫi��7�z,���C-�&̍�oT�a���)��� B"���I�&B\ځ���T|��#�TyK%�JFPs��
3�����n!{z+?í��Iu�Ι��|X���<��M���!�	�۴��w��1S:&!���G���$�Gz;��8� 6<#ܑ�;l��'@��
q��cg���1;A:�n�J��̊���}�خ ��k,�{�X�4��I�>?i�[ly������3y��Q1���4kE�u�Yʑ���$��Z\��5E �ɇ'�)�k�[-Z�(!�ЬL�Qn,�m�ܲv�A���_���y\��fnRF����:�^2X�Hv���.cy���x}��|AB*��N�����31/�ݡ���6B41�1�S���RS"m}�cڠ�XbeJ�d�:��ɚ�V&$���4� !��A��{�A�Tl�������"(��T�&��Q���8�D8�Gw��z�
Ŵ,A�$�R:��@D�m-6�J��T��ibT���I�]b��3�"�?2][^a�
�#Æ���"�����@
̗	�e��K�`��_�u��d!2>�r=*?��ۓWvS")�*]��*��C�cT��3rrh�hd8�df�.!L��,=х>
�I���>=�>I�����
B<d��e���̝��+��] d z�L©{��	���?7�" >bB�.�@E��F��,�,n4���rY��a s���h�*�T���w�B}�~�%�z^;�%���@T�}cS�i��2���oNx��1�����f�(,-I��C���$�~��t���~����D��P�㝎�=L�_�?�qoR&ģ�Y�S���S��̹�-�^����{k���g��烀�	CD�}.��d�k-q-���̖��lt�b6}y�<��#���J�.��F�¹	���` 1����4��aqf5A�>2��4�C\7�3tp"#*�6.4�-f#��1�ׅ�j���	����S�¿a��$'pWV\ �S�cV�x6]F9$�����q?��������hb��s��:��d���=����!��wy��7�+@����\��=$=�(�9N>��?�e����a9Я�Ͻ��Xu�h�WCnd9O�֍�µ2@@&_���7��$�|a��vT���
�^"�����4��$�-��h����x���&*��W�&P"����c�w�o�v������Y|��(�b�7��6Z�,���b{Y%�OY~�D��{)��E�U�A&ٟa����H׊�+*40)�"�Jk��k_gM�O<�qkȵ,g:_�@��;9��t&��G��n�ʛ�$ىN�ѨA�L��a:� 1'^�7����7�0c�3|��}��f���O��k�{�?��ڂ�l���^A�:4{·��D=1��݃[��Mz�,�x�\*F�O�^/���	�Wj� �↪q޵�)� %��^�D̿�w�޶��t�!/ź�}�t�Д*w3����0,�X�a���g�j�6g�D���ϟ�s���Y"Ok�'-σ`n�WF?W8^�q�C�5Ւ�]ۀ1Q�.r����F��!3��^��6˃��6�����k��o�lZ�A���WX"0�x���h��#٣�E�]��+�\NUa?U˥�j�Ŕ��D�wn-�K�$`��Ti��L-
����ihX(��P	�\��-\#�}i���Xb�pX�)���d��$�@:�3Q���9��v0x�b�Q�qL�����x���}�G���.Ie�,���L�	b4Y�̑!֐��"�:\N�5I����B.7�h��Q�@�yLB[����4�2�2�3n�8��d�)S�ӑ�I#i�F��-��~���/ɏK�s��Ig���7���׼	��E��i4����Q�[���e��!O�M:��pt��a�vVt��ͼeU��6�P�h���������J������"��@��r&�"�X�0��Sn2xHAO#i	�(ru%u:wu��<�>&"j�\�loG�ϟ���������W8����o���K�v�Uq���ʎj�3B�uE���������E�%�����-�5�D��JR�Yo�`��D�����bI��c���\��sڞ���7�})+�7��֚!������t������'^�S�dM2)7ιB$lxH�sN��F&��DT��xF��\�Y����Y8�(Y��T�d
�[�7S�4�tњ�s�}��i������F�g��ȣ�nWˋ3냿|j�]���V"�`-sq*:u�\*h*l�>~i��93�go�nn2��#L�Eo;9���^��$�o��(��z�^1o?|�B�B�S����dr�f��"L6�n}�B��y�
�A�>�YVd8@�W�s���W!�L����9j��j]�!+��/ [�p�]
!�
	`�'���z뭴\q�-�Ў�l&Y'��LL�B��%�V�	�ܹA	I���o��o���͉�-A�N��Du,�҂��*�!V��7J�Iʻ;�
���f&��:0�����:��[��r�ݡ��AR�`5B�@2X�w6�Aj@]�Pp�A��E�����B�@���{/e�Y��{�!ϳ\����X>��-G��"��R�� �i��RH�͏���LˉW�`sS�b�O���Hmv	|���z�<��JhZxȀ��c�I���@��X�UH��{H����>�ҡ��<��`2�mR#��i�-�of���,Pq�; %g�"Ac����Y��|_��5�-�d1�|B��"�B�X��E�;ї4)2���!%����a� Z� �8w����@���(��k�r���Mȿ���u1��R0������\@�I48/���/Q�\�}�_A���&J_`-��M����ĥ�~����� H�B�x�~��i���n����B�J.ER<��&�_1y,�~�}@�� �bї��:`������|:����6��P��S�ǂ�]_	����Ѻ��;�\2�߷o�����!�F��}ރeB<Z�U�Kɳ�[d���U�ti����r�CL�*p���x��xH���L7���V@��4�$����nr�x���B�������\^7� ���R��]O ?R�{I�邁[���ظ�$#���_	����k'--\�rb�`���5�@�FYUC<�`J�-�����I�7i�r}i�19�p�s`!����g&�k�ϊ��5`��͖�܈�uiI"(C9��b�^4L��Lb�d�Bư(�ii yU�
������X�𘁔=�``�B��TK��+I��L-�o0~��}�����빦�������@]=�炚�8 ��I�� ����F�G\� A�TGW_v>�Z� �����U^����]jl\�x=,���5����1b�D��3�zC�C�=��~�@�W�e�B�\b_�,5&�&Q��@PBT���pǼ@�	�m�b���!.��5Dp��0�G��e�B#u�}�=���B�.[P��-,�S��O�Rc�M�ףn�U^N�,˻�_G�ռ=�BB~Lj8��y\7�	I$�ϋ}�/��v881��PcktU�ˠN^
z�oB�l��t~X�R��$p4�q�h���p��nVTLn�wz%-�m5
��ur4��*�`^��DH�0Wq��)�p=�$��>B�1��U�5���P�UB�I��xP͓R����LC%�J���'��/���"��aB5OJ��?T�
V    IEND�B`�PK 
     Y�#\rB�. .                  cirkitFile.jsonPK 
     Y�#\                        [ jsons/PK 
     Y�#\Y��c|7  |7                jsons/user_defined.jsonPK 
     Y�#\                        0G images/PK 
     Y�#\��9�� �� /             UG images/04079d65-5a5d-4b08-9f2d-4934008ae210.pngPK 
     Y�#\��ZO%u  %u  /             2+ images/c73ef27d-6394-4828-a75f-205a980bbd83.pngPK 
     Y�#\1�9�c  c  /             �� images/c3d75dd9-81e0-4ecb-9109-310dbcf70c9d.pngPK 
     Y�#\�Q��"  "  /             T� images/c7f8a6b2-5f4f-47a7-84b3-7bbc451b7ab1.pngPK 
     Y�#\q�,��  �  /             ý images/be1ff175-690b-4799-aad0-0ab57f9a01ac.pngPK 
     Y�#\�Vw�    /             �� images/a7a20d0b-f771-49dd-a52a-92c84cdc73c6.pngPK 
     Y�#\�� <   <  /             \� images/e7e47810-abf9-4bb0-84d9-bf12c3babd78.pngPK 
     Y�#\
�  �  /             �	 images/9eaf56c3-a2ed-4703-8e91-9b98c221ec28.pngPK 
     Y�#\VX��<,  <,  /             �) images/5ccbe72c-6fd5-45d2-8118-bee80363f106.pngPK 
     Y�#\��s��  �  /             #V images/e4bf1f14-66df-463a-8792-8567b691137d.pngPK 
     Y�#\q���W W /             )Z images/7c9bed20-c7d7-43dc-b689-820375f46db8.pngPK 
     Y�#\$�3  3  /             �� images/7ade412b-fa94-47ea-987a-d6c9baa14438.pngPK      G  �   